module f_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [13:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'd0: dout <= -'sd587;
        'd1: dout <= 'sd1620;
        'd2: dout <= 'sd1846;
        'd3: dout <= -'sd504;
        'd4: dout <= 'sd213;
        'd5: dout <= 'sd1460;
        'd6: dout <= -'sd771;
        'd7: dout <= -'sd1404;
        'd8: dout <= 'sd711;
        'd9: dout <= -'sd698;
        'd10: dout <= 'sd14;
        'd11: dout <= 'sd923;
        'd12: dout <= -'sd1469;
        'd13: dout <= -'sd2130;
        'd14: dout <= 'sd2097;
        'd15: dout <= -'sd606;
        'd16: dout <= -'sd1346;
        'd17: dout <= 'sd334;
        'd18: dout <= 'sd1357;
        'd19: dout <= -'sd1700;
        'd20: dout <= 'sd2004;
        'd21: dout <= 'sd139;
        'd22: dout <= -'sd415;
        'd23: dout <= -'sd699;
        'd24: dout <= 'sd2171;
        'd25: dout <= -'sd787;
        'd26: dout <= -'sd157;
        'd27: dout <= 'sd1864;
        'd28: dout <= 'sd756;
        'd29: dout <= -'sd665;
        'd30: dout <= 'sd929;
        'd31: dout <= -'sd750;
        'd32: dout <= -'sd2201;
        'd33: dout <= -'sd675;
        'd34: dout <= -'sd1231;
        'd35: dout <= -'sd80;
        'd36: dout <= -'sd138;
        'd37: dout <= -'sd1132;
        'd38: dout <= 'sd957;
        'd39: dout <= 'sd627;
        'd40: dout <= 'sd1125;
        'd41: dout <= -'sd385;
        'd42: dout <= 'sd2263;
        'd43: dout <= -'sd147;
        'd44: dout <= -'sd1257;
        'd45: dout <= -'sd1415;
        'd46: dout <= 'sd622;
        'd47: dout <= 'sd1415;
        'd48: dout <= 'sd1729;
        'd49: dout <= 'sd421;
        'd50: dout <= 'sd1865;
        'd51: dout <= 'sd1529;
        'd52: dout <= 'sd799;
        'd53: dout <= -'sd1637;
        'd54: dout <= -'sd178;
        'd55: dout <= -'sd627;
        'd56: dout <= 'sd1651;
        'd57: dout <= -'sd829;
        'd58: dout <= 'sd1182;
        'd59: dout <= 'sd197;
        'd60: dout <= -'sd1320;
        'd61: dout <= -'sd1533;
        'd62: dout <= 'sd1840;
        'd63: dout <= -'sd1696;
        'd64: dout <= 'sd31;
        'd65: dout <= -'sd1413;
        'd66: dout <= 'sd333;
        'd67: dout <= 'sd29;
        'd68: dout <= -'sd1181;
        'd69: dout <= 'sd1662;
        'd70: dout <= -'sd92;
        'd71: dout <= 'sd1937;
        'd72: dout <= -'sd2164;
        'd73: dout <= 'sd597;
        'd74: dout <= -'sd1997;
        'd75: dout <= -'sd786;
        'd76: dout <= -'sd1438;
        'd77: dout <= 'sd227;
        'd78: dout <= -'sd1475;
        'd79: dout <= 'sd456;
        'd80: dout <= 'sd1907;
        'd81: dout <= 'sd302;
        'd82: dout <= 'sd448;
        'd83: dout <= -'sd32;
        'd84: dout <= 'sd1486;
        'd85: dout <= 'sd2058;
        'd86: dout <= 'sd1235;
        'd87: dout <= 'sd376;
        'd88: dout <= 'sd1600;
        'd89: dout <= 'sd2061;
        'd90: dout <= 'sd1302;
        'd91: dout <= 'sd723;
        'd92: dout <= 'sd801;
        'd93: dout <= -'sd903;
        'd94: dout <= 'sd258;
        'd95: dout <= 'sd1660;
        'd96: dout <= 'sd1715;
        'd97: dout <= -'sd1178;
        'd98: dout <= -'sd1838;
        'd99: dout <= 'sd40;
        'd100: dout <= 'sd1760;
        'd101: dout <= -'sd1884;
        'd102: dout <= 'sd409;
        'd103: dout <= 'sd1385;
        'd104: dout <= -'sd1546;
        'd105: dout <= -'sd694;
        'd106: dout <= -'sd21;
        'd107: dout <= 'sd2292;
        'd108: dout <= 'sd1265;
        'd109: dout <= -'sd168;
        'd110: dout <= 'sd407;
        'd111: dout <= 'sd991;
        'd112: dout <= 'sd519;
        'd113: dout <= -'sd63;
        'd114: dout <= 'sd2182;
        'd115: dout <= -'sd1271;
        'd116: dout <= 'sd1882;
        'd117: dout <= 'sd1414;
        'd118: dout <= 'sd1204;
        'd119: dout <= 'sd374;
        'd120: dout <= -'sd565;
        'd121: dout <= 'sd1387;
        'd122: dout <= 'sd653;
        'd123: dout <= 'sd1978;
        'd124: dout <= 'sd2077;
        'd125: dout <= -'sd853;
        'd126: dout <= 'sd1796;
        'd127: dout <= -'sd977;
        'd128: dout <= -'sd27;
        'd129: dout <= -'sd101;
        'd130: dout <= 'sd1912;
        'd131: dout <= -'sd987;
        'd132: dout <= -'sd174;
        'd133: dout <= 'sd746;
        'd134: dout <= -'sd302;
        'd135: dout <= -'sd2039;
        'd136: dout <= 'sd976;
        'd137: dout <= -'sd749;
        'd138: dout <= 'sd2089;
        'd139: dout <= 'sd555;
        'd140: dout <= 'sd9;
        'd141: dout <= 'sd1368;
        'd142: dout <= 'sd1950;
        'd143: dout <= -'sd187;
        'd144: dout <= -'sd2038;
        'd145: dout <= -'sd863;
        'd146: dout <= 'sd1622;
        'd147: dout <= 'sd572;
        'd148: dout <= -'sd329;
        'd149: dout <= 'sd2026;
        'd150: dout <= -'sd904;
        'd151: dout <= -'sd1897;
        'd152: dout <= 'sd1875;
        'd153: dout <= 'sd1080;
        'd154: dout <= -'sd141;
        'd155: dout <= -'sd1710;
        'd156: dout <= 'sd2143;
        'd157: dout <= -'sd1043;
        'd158: dout <= 'sd1010;
        'd159: dout <= 'sd2021;
        'd160: dout <= -'sd195;
        'd161: dout <= 'sd1113;
        'd162: dout <= 'sd763;
        'd163: dout <= -'sd13;
        'd164: dout <= -'sd215;
        'd165: dout <= -'sd996;
        'd166: dout <= 'sd344;
        'd167: dout <= -'sd842;
        'd168: dout <= 'sd1884;
        'd169: dout <= -'sd1293;
        'd170: dout <= -'sd2277;
        'd171: dout <= -'sd1038;
        'd172: dout <= 'sd1839;
        'd173: dout <= -'sd1737;
        'd174: dout <= 'sd1590;
        'd175: dout <= 'sd64;
        'd176: dout <= -'sd953;
        'd177: dout <= -'sd1413;
        'd178: dout <= -'sd1581;
        'd179: dout <= 'sd378;
        'd180: dout <= 'sd999;
        'd181: dout <= -'sd1544;
        'd182: dout <= 'sd1285;
        'd183: dout <= 'sd138;
        'd184: dout <= 'sd1865;
        'd185: dout <= 'sd541;
        'd186: dout <= 'sd1768;
        'd187: dout <= -'sd1626;
        'd188: dout <= 'sd1742;
        'd189: dout <= 'sd100;
        'd190: dout <= -'sd2005;
        'd191: dout <= 'sd1475;
        'd192: dout <= 'sd1643;
        'd193: dout <= -'sd360;
        'd194: dout <= -'sd1697;
        'd195: dout <= -'sd894;
        'd196: dout <= -'sd1976;
        'd197: dout <= -'sd2045;
        'd198: dout <= 'sd1801;
        'd199: dout <= -'sd1017;
        'd200: dout <= 'sd212;
        'd201: dout <= 'sd1831;
        'd202: dout <= -'sd1437;
        'd203: dout <= -'sd556;
        'd204: dout <= 'sd1447;
        'd205: dout <= -'sd1697;
        'd206: dout <= -'sd332;
        'd207: dout <= -'sd1058;
        'd208: dout <= -'sd2214;
        'd209: dout <= 'sd2295;
        'd210: dout <= -'sd961;
        'd211: dout <= -'sd80;
        'd212: dout <= 'sd1703;
        'd213: dout <= 'sd1817;
        'd214: dout <= -'sd1272;
        'd215: dout <= 'sd904;
        'd216: dout <= 'sd1100;
        'd217: dout <= -'sd1959;
        'd218: dout <= 'sd507;
        'd219: dout <= 'sd1452;
        'd220: dout <= -'sd1107;
        'd221: dout <= -'sd1909;
        'd222: dout <= -'sd814;
        'd223: dout <= 'sd552;
        'd224: dout <= 'sd1469;
        'd225: dout <= 'sd1813;
        'd226: dout <= 'sd1316;
        'd227: dout <= -'sd24;
        'd228: dout <= -'sd93;
        'd229: dout <= 'sd1110;
        'd230: dout <= 'sd1328;
        'd231: dout <= 'sd2031;
        'd232: dout <= 'sd1385;
        'd233: dout <= -'sd735;
        'd234: dout <= 'sd2168;
        'd235: dout <= -'sd1936;
        'd236: dout <= -'sd1245;
        'd237: dout <= 'sd709;
        'd238: dout <= -'sd1346;
        'd239: dout <= -'sd838;
        'd240: dout <= -'sd350;
        'd241: dout <= 'sd1542;
        'd242: dout <= -'sd177;
        'd243: dout <= -'sd2113;
        'd244: dout <= -'sd1077;
        'd245: dout <= -'sd1018;
        'd246: dout <= -'sd308;
        'd247: dout <= -'sd693;
        'd248: dout <= -'sd1923;
        'd249: dout <= -'sd483;
        'd250: dout <= -'sd1446;
        'd251: dout <= 'sd1084;
        'd252: dout <= 'sd1861;
        'd253: dout <= -'sd1502;
        'd254: dout <= 'sd1210;
        'd255: dout <= -'sd494;
        'd256: dout <= -'sd339;
        'd257: dout <= -'sd6;
        'd258: dout <= 'sd1000;
        'd259: dout <= 'sd557;
        'd260: dout <= 'sd603;
        'd261: dout <= 'sd514;
        'd262: dout <= -'sd1886;
        'd263: dout <= 'sd1199;
        'd264: dout <= -'sd1023;
        'd265: dout <= -'sd1717;
        'd266: dout <= 'sd37;
        'd267: dout <= 'sd582;
        'd268: dout <= -'sd1279;
        'd269: dout <= 'sd1463;
        'd270: dout <= -'sd1487;
        'd271: dout <= -'sd1251;
        'd272: dout <= -'sd892;
        'd273: dout <= 'sd490;
        'd274: dout <= -'sd687;
        'd275: dout <= -'sd379;
        'd276: dout <= 'sd397;
        'd277: dout <= 'sd662;
        'd278: dout <= -'sd783;
        'd279: dout <= -'sd1485;
        'd280: dout <= 'sd868;
        'd281: dout <= 'sd246;
        'd282: dout <= 'sd1341;
        'd283: dout <= -'sd2060;
        'd284: dout <= 'sd239;
        'd285: dout <= 'sd1104;
        'd286: dout <= 'sd790;
        'd287: dout <= -'sd151;
        'd288: dout <= -'sd420;
        'd289: dout <= -'sd929;
        'd290: dout <= 'sd327;
        'd291: dout <= -'sd1381;
        'd292: dout <= 'sd599;
        'd293: dout <= -'sd1152;
        'd294: dout <= -'sd1538;
        'd295: dout <= 'sd671;
        'd296: dout <= 'sd1443;
        'd297: dout <= -'sd884;
        'd298: dout <= 'sd168;
        'd299: dout <= -'sd741;
        'd300: dout <= -'sd590;
        'd301: dout <= 'sd1362;
        'd302: dout <= -'sd1101;
        'd303: dout <= 'sd750;
        'd304: dout <= -'sd311;
        'd305: dout <= 'sd565;
        'd306: dout <= 'sd2150;
        'd307: dout <= 'sd63;
        'd308: dout <= -'sd961;
        'd309: dout <= 'sd608;
        'd310: dout <= 'sd1919;
        'd311: dout <= -'sd79;
        'd312: dout <= -'sd870;
        'd313: dout <= 'sd1648;
        'd314: dout <= 'sd477;
        'd315: dout <= 'sd1792;
        'd316: dout <= 'sd54;
        'd317: dout <= -'sd944;
        'd318: dout <= -'sd1856;
        'd319: dout <= 'sd230;
        'd320: dout <= -'sd1419;
        'd321: dout <= -'sd401;
        'd322: dout <= -'sd2238;
        'd323: dout <= 'sd520;
        'd324: dout <= -'sd24;
        'd325: dout <= 'sd713;
        'd326: dout <= 'sd2220;
        'd327: dout <= 'sd903;
        'd328: dout <= -'sd1849;
        'd329: dout <= -'sd1893;
        'd330: dout <= 'sd765;
        'd331: dout <= -'sd382;
        'd332: dout <= -'sd665;
        'd333: dout <= -'sd81;
        'd334: dout <= 'sd1865;
        'd335: dout <= -'sd1640;
        'd336: dout <= -'sd508;
        'd337: dout <= -'sd1928;
        'd338: dout <= 'sd1692;
        'd339: dout <= -'sd2045;
        'd340: dout <= 'sd450;
        'd341: dout <= 'sd1321;
        'd342: dout <= -'sd1068;
        'd343: dout <= -'sd336;
        'd344: dout <= 'sd855;
        'd345: dout <= 'sd2270;
        'd346: dout <= 'sd1293;
        'd347: dout <= 'sd2244;
        'd348: dout <= -'sd554;
        'd349: dout <= 'sd1325;
        'd350: dout <= -'sd783;
        'd351: dout <= 'sd1357;
        'd352: dout <= -'sd297;
        'd353: dout <= -'sd1883;
        'd354: dout <= -'sd767;
        'd355: dout <= -'sd1937;
        'd356: dout <= 'sd1664;
        'd357: dout <= 'sd214;
        'd358: dout <= 'sd1434;
        'd359: dout <= 'sd1452;
        'd360: dout <= -'sd770;
        'd361: dout <= 'sd1162;
        'd362: dout <= 'sd1078;
        'd363: dout <= 'sd1665;
        'd364: dout <= 'sd2241;
        'd365: dout <= -'sd124;
        'd366: dout <= -'sd1698;
        'd367: dout <= 'sd2035;
        'd368: dout <= 'sd1863;
        'd369: dout <= -'sd2243;
        'd370: dout <= 'sd2291;
        'd371: dout <= -'sd1580;
        'd372: dout <= 'sd1179;
        'd373: dout <= 'sd1419;
        'd374: dout <= -'sd1099;
        'd375: dout <= -'sd1364;
        'd376: dout <= 'sd1048;
        'd377: dout <= 'sd1203;
        'd378: dout <= -'sd51;
        'd379: dout <= -'sd1306;
        'd380: dout <= -'sd2265;
        'd381: dout <= 'sd2003;
        'd382: dout <= -'sd420;
        'd383: dout <= 'sd1871;
        'd384: dout <= 'sd618;
        'd385: dout <= 'sd2048;
        'd386: dout <= 'sd2173;
        'd387: dout <= 'sd1591;
        'd388: dout <= -'sd1319;
        'd389: dout <= 'sd588;
        'd390: dout <= -'sd345;
        'd391: dout <= -'sd18;
        'd392: dout <= -'sd795;
        'd393: dout <= -'sd357;
        'd394: dout <= -'sd880;
        'd395: dout <= 'sd1678;
        'd396: dout <= 'sd84;
        'd397: dout <= 'sd752;
        'd398: dout <= 'sd680;
        'd399: dout <= 'sd1333;
        'd400: dout <= 'sd1174;
        'd401: dout <= 'sd1728;
        'd402: dout <= -'sd476;
        'd403: dout <= -'sd1788;
        'd404: dout <= 'sd1840;
        'd405: dout <= -'sd789;
        'd406: dout <= 'sd1677;
        'd407: dout <= 'sd496;
        'd408: dout <= -'sd407;
        'd409: dout <= 'sd320;
        'd410: dout <= 'sd1643;
        'd411: dout <= 'sd2068;
        'd412: dout <= 'sd321;
        'd413: dout <= 'sd1543;
        'd414: dout <= 'sd98;
        'd415: dout <= -'sd832;
        'd416: dout <= -'sd278;
        'd417: dout <= -'sd2168;
        'd418: dout <= -'sd296;
        'd419: dout <= 'sd981;
        'd420: dout <= -'sd922;
        'd421: dout <= 'sd179;
        'd422: dout <= -'sd1691;
        'd423: dout <= 'sd2011;
        'd424: dout <= 'sd1512;
        'd425: dout <= 'sd1774;
        'd426: dout <= -'sd2017;
        'd427: dout <= -'sd2274;
        'd428: dout <= 'sd1428;
        'd429: dout <= -'sd1303;
        'd430: dout <= -'sd121;
        'd431: dout <= -'sd365;
        'd432: dout <= 'sd993;
        'd433: dout <= -'sd1003;
        'd434: dout <= 'sd1140;
        'd435: dout <= 'sd330;
        'd436: dout <= 'sd1739;
        'd437: dout <= 'sd559;
        'd438: dout <= -'sd1801;
        'd439: dout <= 'sd68;
        'd440: dout <= 'sd902;
        'd441: dout <= 'sd1947;
        'd442: dout <= -'sd1265;
        'd443: dout <= -'sd1681;
        'd444: dout <= 'sd2158;
        'd445: dout <= 'sd652;
        'd446: dout <= 'sd464;
        'd447: dout <= 'sd740;
        'd448: dout <= -'sd384;
        'd449: dout <= 'sd534;
        'd450: dout <= -'sd853;
        'd451: dout <= -'sd555;
        'd452: dout <= -'sd249;
        'd453: dout <= 'sd441;
        'd454: dout <= 'sd989;
        'd455: dout <= 'sd173;
        'd456: dout <= 'sd1984;
        'd457: dout <= 'sd797;
        'd458: dout <= 'sd1006;
        'd459: dout <= -'sd176;
        'd460: dout <= 'sd1607;
        'd461: dout <= 'sd417;
        'd462: dout <= -'sd956;
        'd463: dout <= 'sd334;
        'd464: dout <= -'sd2056;
        'd465: dout <= -'sd634;
        'd466: dout <= 'sd1067;
        'd467: dout <= 'sd131;
        'd468: dout <= -'sd1958;
        'd469: dout <= -'sd1480;
        'd470: dout <= -'sd2028;
        'd471: dout <= 'sd1073;
        'd472: dout <= -'sd313;
        'd473: dout <= -'sd1894;
        'd474: dout <= -'sd560;
        'd475: dout <= 'sd2202;
        'd476: dout <= 'sd415;
        'd477: dout <= -'sd1332;
        'd478: dout <= -'sd53;
        'd479: dout <= -'sd340;
        'd480: dout <= 'sd1437;
        'd481: dout <= 'sd1711;
        'd482: dout <= 'sd1863;
        'd483: dout <= -'sd1560;
        'd484: dout <= 'sd404;
        'd485: dout <= 'sd1240;
        'd486: dout <= -'sd977;
        'd487: dout <= 'sd774;
        'd488: dout <= 'sd1423;
        'd489: dout <= 'sd716;
        'd490: dout <= -'sd1573;
        'd491: dout <= -'sd2146;
        'd492: dout <= 'sd393;
        'd493: dout <= -'sd1457;
        'd494: dout <= -'sd2165;
        'd495: dout <= -'sd1956;
        'd496: dout <= -'sd1438;
        'd497: dout <= 'sd1565;
        'd498: dout <= 'sd1365;
        'd499: dout <= 'sd1968;
        'd500: dout <= -'sd814;
        'd501: dout <= -'sd956;
        'd502: dout <= -'sd1120;
        'd503: dout <= 'sd1143;
        'd504: dout <= -'sd224;
        'd505: dout <= -'sd1600;
        'd506: dout <= -'sd2194;
        'd507: dout <= -'sd800;
        'd508: dout <= 'sd689;
        'd509: dout <= 'sd1265;
        'd510: dout <= -'sd1366;
        'd511: dout <= 'sd1545;
        'd512: dout <= 'sd1305;
        'd513: dout <= 'sd1331;
        'd514: dout <= -'sd27;
        'd515: dout <= -'sd952;
        'd516: dout <= -'sd812;
        'd517: dout <= -'sd1821;
        'd518: dout <= -'sd1767;
        'd519: dout <= 'sd959;
        'd520: dout <= 'sd1551;
        'd521: dout <= -'sd2139;
        'd522: dout <= -'sd701;
        'd523: dout <= 'sd503;
        'd524: dout <= -'sd1947;
        'd525: dout <= -'sd410;
        'd526: dout <= -'sd479;
        'd527: dout <= 'sd633;
        'd528: dout <= 'sd1930;
        'd529: dout <= 'sd1338;
        'd530: dout <= -'sd1393;
        'd531: dout <= -'sd1504;
        'd532: dout <= 'sd1378;
        'd533: dout <= -'sd1365;
        'd534: dout <= -'sd939;
        'd535: dout <= 'sd1827;
        'd536: dout <= 'sd1471;
        'd537: dout <= -'sd1982;
        'd538: dout <= 'sd784;
        'd539: dout <= 'sd1083;
        'd540: dout <= 'sd524;
        'd541: dout <= 'sd1896;
        'd542: dout <= 'sd302;
        'd543: dout <= 'sd136;
        'd544: dout <= -'sd887;
        'd545: dout <= 'sd476;
        'd546: dout <= 'sd1245;
        'd547: dout <= 'sd1776;
        'd548: dout <= -'sd1813;
        'd549: dout <= -'sd1427;
        'd550: dout <= -'sd36;
        'd551: dout <= 'sd1837;
        'd552: dout <= -'sd1805;
        'd553: dout <= -'sd1607;
        'd554: dout <= -'sd1772;
        'd555: dout <= -'sd680;
        'd556: dout <= -'sd364;
        'd557: dout <= 'sd1171;
        'd558: dout <= -'sd678;
        'd559: dout <= -'sd890;
        'd560: dout <= -'sd1402;
        'd561: dout <= -'sd280;
        'd562: dout <= -'sd174;
        'd563: dout <= 'sd915;
        'd564: dout <= 'sd1797;
        'd565: dout <= 'sd1313;
        'd566: dout <= -'sd820;
        'd567: dout <= 'sd229;
        'd568: dout <= 'sd1850;
        'd569: dout <= 'sd1137;
        'd570: dout <= 'sd294;
        'd571: dout <= -'sd1274;
        'd572: dout <= 'sd1386;
        'd573: dout <= -'sd2146;
        'd574: dout <= 'sd1226;
        'd575: dout <= -'sd303;
        'd576: dout <= 'sd1721;
        'd577: dout <= 'sd2109;
        'd578: dout <= 'sd2064;
        'd579: dout <= 'sd956;
        'd580: dout <= -'sd195;
        'd581: dout <= 'sd663;
        'd582: dout <= 'sd1840;
        'd583: dout <= 'sd1820;
        'd584: dout <= 'sd882;
        'd585: dout <= -'sd1522;
        'd586: dout <= 'sd1217;
        'd587: dout <= -'sd1043;
        'd588: dout <= -'sd591;
        'd589: dout <= -'sd1440;
        'd590: dout <= 'sd515;
        'd591: dout <= 'sd1657;
        'd592: dout <= 'sd818;
        'd593: dout <= -'sd1893;
        'd594: dout <= -'sd1339;
        'd595: dout <= 'sd2056;
        'd596: dout <= 'sd1237;
        'd597: dout <= 'sd1688;
        'd598: dout <= -'sd1203;
        'd599: dout <= 'sd1830;
        'd600: dout <= -'sd707;
        'd601: dout <= 'sd720;
        'd602: dout <= -'sd1351;
        'd603: dout <= -'sd1268;
        'd604: dout <= -'sd221;
        'd605: dout <= 'sd1986;
        'd606: dout <= -'sd2024;
        'd607: dout <= 'sd1271;
        'd608: dout <= -'sd1683;
        'd609: dout <= 'sd1242;
        'd610: dout <= -'sd1949;
        'd611: dout <= -'sd2244;
        'd612: dout <= -'sd2210;
        'd613: dout <= 'sd1748;
        'd614: dout <= 'sd420;
        'd615: dout <= 'sd537;
        'd616: dout <= 'sd1737;
        'd617: dout <= 'sd1746;
        'd618: dout <= -'sd1687;
        'd619: dout <= -'sd1259;
        'd620: dout <= 'sd972;
        'd621: dout <= -'sd614;
        'd622: dout <= 'sd2102;
        'd623: dout <= 'sd1672;
        'd624: dout <= -'sd1212;
        'd625: dout <= 'sd1011;
        'd626: dout <= 'sd823;
        'd627: dout <= -'sd639;
        'd628: dout <= 'sd2274;
        'd629: dout <= -'sd1577;
        'd630: dout <= 'sd1530;
        'd631: dout <= 'sd241;
        'd632: dout <= -'sd773;
        'd633: dout <= -'sd616;
        'd634: dout <= -'sd759;
        'd635: dout <= -'sd410;
        'd636: dout <= -'sd1653;
        'd637: dout <= 'sd787;
        'd638: dout <= -'sd1558;
        'd639: dout <= 'sd2184;
        'd640: dout <= -'sd1723;
        'd641: dout <= 'sd311;
        'd642: dout <= -'sd486;
        'd643: dout <= 'sd72;
        'd644: dout <= -'sd1963;
        'd645: dout <= 'sd477;
        'd646: dout <= 'sd2102;
        'd647: dout <= 'sd1388;
        'd648: dout <= -'sd1438;
        'd649: dout <= 'sd2248;
        'd650: dout <= -'sd810;
        'd651: dout <= 'sd1183;
        'd652: dout <= 'sd931;
        'd653: dout <= -'sd820;
        'd654: dout <= 'sd1716;
        'd655: dout <= 'sd1705;
        'd656: dout <= -'sd903;
        'd657: dout <= 'sd2247;
        'd658: dout <= -'sd341;
        'd659: dout <= -'sd1320;
        'd660: dout <= 'sd1568;
        'd661: dout <= 'sd1825;
        'd662: dout <= 'sd961;
        'd663: dout <= -'sd1416;
        'd664: dout <= -'sd1691;
        'd665: dout <= -'sd1627;
        'd666: dout <= 'sd233;
        'd667: dout <= 'sd412;
        'd668: dout <= 'sd1578;
        'd669: dout <= 'sd2026;
        'd670: dout <= -'sd1222;
        'd671: dout <= 'sd934;
        'd672: dout <= 'sd1595;
        'd673: dout <= -'sd810;
        'd674: dout <= -'sd120;
        'd675: dout <= -'sd1590;
        'd676: dout <= -'sd276;
        'd677: dout <= 'sd279;
        'd678: dout <= -'sd904;
        'd679: dout <= -'sd1206;
        'd680: dout <= -'sd475;
        'd681: dout <= -'sd38;
        'd682: dout <= 'sd540;
        'd683: dout <= 'sd1196;
        'd684: dout <= -'sd1998;
        'd685: dout <= 'sd394;
        'd686: dout <= 'sd1690;
        'd687: dout <= -'sd1777;
        'd688: dout <= 'sd2253;
        'd689: dout <= 'sd1890;
        'd690: dout <= -'sd137;
        'd691: dout <= -'sd1969;
        'd692: dout <= 'sd563;
        'd693: dout <= -'sd533;
        'd694: dout <= -'sd563;
        'd695: dout <= 'sd717;
        'd696: dout <= -'sd1696;
        'd697: dout <= 'sd768;
        'd698: dout <= -'sd197;
        'd699: dout <= -'sd1528;
        'd700: dout <= 'sd196;
        'd701: dout <= 'sd1643;
        'd702: dout <= -'sd40;
        'd703: dout <= 'sd1404;
        'd704: dout <= 'sd10;
        'd705: dout <= 'sd2145;
        'd706: dout <= 'sd2052;
        'd707: dout <= 'sd1457;
        'd708: dout <= -'sd1268;
        'd709: dout <= -'sd2232;
        'd710: dout <= -'sd1375;
        'd711: dout <= -'sd1738;
        'd712: dout <= -'sd431;
        'd713: dout <= 'sd410;
        'd714: dout <= -'sd1523;
        'd715: dout <= 'sd871;
        'd716: dout <= -'sd97;
        'd717: dout <= -'sd78;
        'd718: dout <= -'sd375;
        'd719: dout <= -'sd1202;
        'd720: dout <= 'sd1686;
        'd721: dout <= -'sd924;
        'd722: dout <= 'sd2186;
        'd723: dout <= 'sd1339;
        'd724: dout <= -'sd124;
        'd725: dout <= 'sd533;
        'd726: dout <= 'sd121;
        'd727: dout <= -'sd651;
        'd728: dout <= 'sd2128;
        'd729: dout <= 'sd1767;
        'd730: dout <= -'sd2267;
        'd731: dout <= 'sd1954;
        'd732: dout <= 'sd1255;
        'd733: dout <= 'sd618;
        'd734: dout <= 'sd1886;
        'd735: dout <= -'sd423;
        'd736: dout <= -'sd1096;
        'd737: dout <= 'sd1901;
        'd738: dout <= -'sd1584;
        'd739: dout <= -'sd2220;
        'd740: dout <= -'sd1245;
        'd741: dout <= 'sd347;
        'd742: dout <= -'sd759;
        'd743: dout <= 'sd1227;
        'd744: dout <= 'sd117;
        'd745: dout <= 'sd667;
        'd746: dout <= -'sd2119;
        'd747: dout <= -'sd932;
        'd748: dout <= -'sd1802;
        'd749: dout <= 'sd1968;
        'd750: dout <= 'sd1785;
        'd751: dout <= 'sd1779;
        'd752: dout <= 'sd1211;
        'd753: dout <= 'sd1511;
        'd754: dout <= -'sd285;
        'd755: dout <= -'sd1118;
        'd756: dout <= 'sd2122;
        'd757: dout <= 'sd320;
        'd758: dout <= 'sd666;
        'd759: dout <= -'sd1449;
        'd760: dout <= -'sd233;
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module g_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [13:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'd0: dout <= 'sd168;
        'd1: dout <= 'sd97;
        'd2: dout <= 'sd630;
        'd3: dout <= 'sd1025;
        'd4: dout <= 'sd338;
        'd5: dout <= 'sd1322;
        'd6: dout <= -'sd784;
        'd7: dout <= 'sd1242;
        'd8: dout <= 'sd1942;
        'd9: dout <= -'sd1352;
        'd10: dout <= -'sd1444;
        'd11: dout <= 'sd357;
        'd12: dout <= -'sd1331;
        'd13: dout <= -'sd960;
        'd14: dout <= -'sd2210;
        'd15: dout <= 'sd2207;
        'd16: dout <= -'sd390;
        'd17: dout <= -'sd1533;
        'd18: dout <= -'sd1486;
        'd19: dout <= -'sd1778;
        'd20: dout <= -'sd279;
        'd21: dout <= -'sd605;
        'd22: dout <= 'sd1545;
        'd23: dout <= 'sd2177;
        'd24: dout <= -'sd1033;
        'd25: dout <= 'sd1899;
        'd26: dout <= 'sd1405;
        'd27: dout <= -'sd661;
        'd28: dout <= 'sd1014;
        'd29: dout <= 'sd762;
        'd30: dout <= -'sd897;
        'd31: dout <= -'sd568;
        'd32: dout <= 'sd1967;
        'd33: dout <= 'sd733;
        'd34: dout <= -'sd1104;
        'd35: dout <= -'sd129;
        'd36: dout <= -'sd513;
        'd37: dout <= 'sd728;
        'd38: dout <= -'sd769;
        'd39: dout <= 'sd96;
        'd40: dout <= -'sd1390;
        'd41: dout <= -'sd1382;
        'd42: dout <= -'sd35;
        'd43: dout <= 'sd2237;
        'd44: dout <= -'sd1419;
        'd45: dout <= 'sd421;
        'd46: dout <= -'sd1037;
        'd47: dout <= -'sd140;
        'd48: dout <= 'sd793;
        'd49: dout <= -'sd1970;
        'd50: dout <= -'sd1843;
        'd51: dout <= 'sd1899;
        'd52: dout <= 'sd1662;
        'd53: dout <= -'sd1025;
        'd54: dout <= 'sd215;
        'd55: dout <= 'sd1112;
        'd56: dout <= -'sd1812;
        'd57: dout <= -'sd1452;
        'd58: dout <= -'sd43;
        'd59: dout <= 'sd1935;
        'd60: dout <= -'sd411;
        'd61: dout <= 'sd1679;
        'd62: dout <= 'sd859;
        'd63: dout <= 'sd2062;
        'd64: dout <= 'sd1674;
        'd65: dout <= 'sd603;
        'd66: dout <= -'sd1930;
        'd67: dout <= 'sd881;
        'd68: dout <= -'sd428;
        'd69: dout <= -'sd1554;
        'd70: dout <= 'sd797;
        'd71: dout <= -'sd11;
        'd72: dout <= -'sd721;
        'd73: dout <= -'sd2290;
        'd74: dout <= 'sd1678;
        'd75: dout <= -'sd971;
        'd76: dout <= -'sd1305;
        'd77: dout <= 'sd706;
        'd78: dout <= 'sd609;
        'd79: dout <= 'sd1655;
        'd80: dout <= 'sd638;
        'd81: dout <= 'sd1622;
        'd82: dout <= 'sd1364;
        'd83: dout <= 'sd1070;
        'd84: dout <= -'sd2013;
        'd85: dout <= 'sd879;
        'd86: dout <= -'sd1862;
        'd87: dout <= 'sd2195;
        'd88: dout <= 'sd275;
        'd89: dout <= 'sd1826;
        'd90: dout <= 'sd1079;
        'd91: dout <= -'sd183;
        'd92: dout <= 'sd808;
        'd93: dout <= 'sd2268;
        'd94: dout <= -'sd807;
        'd95: dout <= -'sd1373;
        'd96: dout <= 'sd1684;
        'd97: dout <= -'sd286;
        'd98: dout <= 'sd1316;
        'd99: dout <= -'sd2097;
        'd100: dout <= -'sd672;
        'd101: dout <= -'sd1422;
        'd102: dout <= 'sd741;
        'd103: dout <= -'sd1926;
        'd104: dout <= 'sd1696;
        'd105: dout <= -'sd561;
        'd106: dout <= 'sd1576;
        'd107: dout <= -'sd1864;
        'd108: dout <= 'sd1362;
        'd109: dout <= -'sd678;
        'd110: dout <= 'sd97;
        'd111: dout <= -'sd2243;
        'd112: dout <= -'sd1577;
        'd113: dout <= 'sd224;
        'd114: dout <= -'sd751;
        'd115: dout <= -'sd1056;
        'd116: dout <= -'sd1156;
        'd117: dout <= 'sd2266;
        'd118: dout <= 'sd1090;
        'd119: dout <= -'sd1368;
        'd120: dout <= -'sd1578;
        'd121: dout <= -'sd1896;
        'd122: dout <= 'sd2214;
        'd123: dout <= 'sd821;
        'd124: dout <= -'sd1345;
        'd125: dout <= 'sd1486;
        'd126: dout <= 'sd527;
        'd127: dout <= 'sd4;
        'd128: dout <= 'sd2006;
        'd129: dout <= 'sd374;
        'd130: dout <= 'sd240;
        'd131: dout <= 'sd1342;
        'd132: dout <= -'sd701;
        'd133: dout <= 'sd2013;
        'd134: dout <= 'sd934;
        'd135: dout <= 'sd995;
        'd136: dout <= -'sd215;
        'd137: dout <= 'sd1674;
        'd138: dout <= 'sd1119;
        'd139: dout <= 'sd829;
        'd140: dout <= -'sd732;
        'd141: dout <= -'sd868;
        'd142: dout <= -'sd1695;
        'd143: dout <= 'sd998;
        'd144: dout <= -'sd1914;
        'd145: dout <= 'sd1847;
        'd146: dout <= -'sd1077;
        'd147: dout <= -'sd1033;
        'd148: dout <= 'sd963;
        'd149: dout <= -'sd2077;
        'd150: dout <= -'sd1304;
        'd151: dout <= -'sd466;
        'd152: dout <= -'sd2045;
        'd153: dout <= 'sd566;
        'd154: dout <= 'sd197;
        'd155: dout <= -'sd300;
        'd156: dout <= 'sd1984;
        'd157: dout <= -'sd938;
        'd158: dout <= -'sd2129;
        'd159: dout <= 'sd1674;
        'd160: dout <= 'sd214;
        'd161: dout <= -'sd1497;
        'd162: dout <= 'sd1681;
        'd163: dout <= 'sd1484;
        'd164: dout <= 'sd249;
        'd165: dout <= 'sd1195;
        'd166: dout <= -'sd61;
        'd167: dout <= -'sd1784;
        'd168: dout <= 'sd748;
        'd169: dout <= -'sd309;
        'd170: dout <= 'sd1289;
        'd171: dout <= -'sd1978;
        'd172: dout <= 'sd412;
        'd173: dout <= 'sd1546;
        'd174: dout <= -'sd1070;
        'd175: dout <= 'sd1071;
        'd176: dout <= -'sd2103;
        'd177: dout <= -'sd83;
        'd178: dout <= 'sd1420;
        'd179: dout <= 'sd2094;
        'd180: dout <= 'sd2176;
        'd181: dout <= -'sd1590;
        'd182: dout <= 'sd1954;
        'd183: dout <= 'sd76;
        'd184: dout <= 'sd705;
        'd185: dout <= 'sd1263;
        'd186: dout <= 'sd782;
        'd187: dout <= 'sd31;
        'd188: dout <= -'sd239;
        'd189: dout <= -'sd913;
        'd190: dout <= 'sd1662;
        'd191: dout <= -'sd1256;
        'd192: dout <= 'sd1158;
        'd193: dout <= -'sd410;
        'd194: dout <= -'sd2158;
        'd195: dout <= 'sd2050;
        'd196: dout <= 'sd321;
        'd197: dout <= -'sd138;
        'd198: dout <= -'sd2153;
        'd199: dout <= 'sd1798;
        'd200: dout <= 'sd1890;
        'd201: dout <= -'sd2222;
        'd202: dout <= -'sd242;
        'd203: dout <= 'sd1151;
        'd204: dout <= 'sd520;
        'd205: dout <= 'sd1418;
        'd206: dout <= 'sd153;
        'd207: dout <= 'sd773;
        'd208: dout <= 'sd1892;
        'd209: dout <= 'sd1373;
        'd210: dout <= 'sd164;
        'd211: dout <= -'sd326;
        'd212: dout <= -'sd723;
        'd213: dout <= -'sd642;
        'd214: dout <= -'sd1291;
        'd215: dout <= 'sd10;
        'd216: dout <= -'sd2025;
        'd217: dout <= 'sd1440;
        'd218: dout <= 'sd1650;
        'd219: dout <= 'sd874;
        'd220: dout <= 'sd703;
        'd221: dout <= -'sd457;
        'd222: dout <= -'sd1969;
        'd223: dout <= -'sd19;
        'd224: dout <= 'sd2141;
        'd225: dout <= 'sd2131;
        'd226: dout <= -'sd1689;
        'd227: dout <= -'sd1303;
        'd228: dout <= -'sd158;
        'd229: dout <= -'sd1483;
        'd230: dout <= 'sd1399;
        'd231: dout <= -'sd227;
        'd232: dout <= 'sd1223;
        'd233: dout <= 'sd2240;
        'd234: dout <= -'sd1733;
        'd235: dout <= 'sd349;
        'd236: dout <= 'sd1169;
        'd237: dout <= -'sd948;
        'd238: dout <= -'sd1196;
        'd239: dout <= -'sd390;
        'd240: dout <= -'sd274;
        'd241: dout <= -'sd1495;
        'd242: dout <= -'sd1339;
        'd243: dout <= 'sd355;
        'd244: dout <= -'sd1431;
        'd245: dout <= 'sd443;
        'd246: dout <= -'sd1510;
        'd247: dout <= -'sd1019;
        'd248: dout <= 'sd1863;
        'd249: dout <= -'sd1360;
        'd250: dout <= 'sd1622;
        'd251: dout <= 'sd1532;
        'd252: dout <= 'sd1384;
        'd253: dout <= -'sd1292;
        'd254: dout <= 'sd1246;
        'd255: dout <= 'sd952;
        'd256: dout <= 'sd117;
        'd257: dout <= 'sd395;
        'd258: dout <= -'sd516;
        'd259: dout <= -'sd1458;
        'd260: dout <= -'sd682;
        'd261: dout <= -'sd2204;
        'd262: dout <= 'sd674;
        'd263: dout <= 'sd331;
        'd264: dout <= -'sd1960;
        'd265: dout <= 'sd1400;
        'd266: dout <= 'sd254;
        'd267: dout <= 'sd1904;
        'd268: dout <= 'sd1039;
        'd269: dout <= -'sd1052;
        'd270: dout <= 'sd269;
        'd271: dout <= 'sd1786;
        'd272: dout <= 'sd1680;
        'd273: dout <= 'sd74;
        'd274: dout <= -'sd618;
        'd275: dout <= -'sd1487;
        'd276: dout <= 'sd316;
        'd277: dout <= 'sd1265;
        'd278: dout <= -'sd1795;
        'd279: dout <= 'sd1424;
        'd280: dout <= -'sd1805;
        'd281: dout <= -'sd1889;
        'd282: dout <= 'sd481;
        'd283: dout <= -'sd309;
        'd284: dout <= 'sd1830;
        'd285: dout <= 'sd69;
        'd286: dout <= -'sd2196;
        'd287: dout <= -'sd276;
        'd288: dout <= -'sd1816;
        'd289: dout <= 'sd1853;
        'd290: dout <= 'sd2275;
        'd291: dout <= -'sd722;
        'd292: dout <= -'sd393;
        'd293: dout <= 'sd320;
        'd294: dout <= -'sd325;
        'd295: dout <= -'sd552;
        'd296: dout <= 'sd742;
        'd297: dout <= -'sd294;
        'd298: dout <= 'sd2119;
        'd299: dout <= -'sd1287;
        'd300: dout <= 'sd879;
        'd301: dout <= 'sd1672;
        'd302: dout <= -'sd2044;
        'd303: dout <= 'sd1684;
        'd304: dout <= 'sd2069;
        'd305: dout <= 'sd1548;
        'd306: dout <= -'sd1529;
        'd307: dout <= 'sd43;
        'd308: dout <= -'sd2061;
        'd309: dout <= -'sd2052;
        'd310: dout <= 'sd1451;
        'd311: dout <= 'sd140;
        'd312: dout <= 'sd1895;
        'd313: dout <= -'sd2130;
        'd314: dout <= 'sd2286;
        'd315: dout <= -'sd1892;
        'd316: dout <= 'sd216;
        'd317: dout <= 'sd1412;
        'd318: dout <= 'sd1622;
        'd319: dout <= 'sd1672;
        'd320: dout <= 'sd245;
        'd321: dout <= 'sd448;
        'd322: dout <= -'sd706;
        'd323: dout <= -'sd850;
        'd324: dout <= -'sd932;
        'd325: dout <= -'sd179;
        'd326: dout <= 'sd771;
        'd327: dout <= -'sd2235;
        'd328: dout <= -'sd1622;
        'd329: dout <= 'sd271;
        'd330: dout <= -'sd1290;
        'd331: dout <= 'sd392;
        'd332: dout <= 'sd22;
        'd333: dout <= -'sd1649;
        'd334: dout <= 'sd1727;
        'd335: dout <= -'sd833;
        'd336: dout <= -'sd1742;
        'd337: dout <= -'sd1328;
        'd338: dout <= 'sd1463;
        'd339: dout <= 'sd1864;
        'd340: dout <= -'sd557;
        'd341: dout <= -'sd1643;
        'd342: dout <= -'sd1652;
        'd343: dout <= -'sd592;
        'd344: dout <= 'sd125;
        'd345: dout <= 'sd1816;
        'd346: dout <= 'sd1628;
        'd347: dout <= -'sd1668;
        'd348: dout <= -'sd574;
        'd349: dout <= -'sd1996;
        'd350: dout <= 'sd143;
        'd351: dout <= -'sd2103;
        'd352: dout <= 'sd2022;
        'd353: dout <= 'sd2143;
        'd354: dout <= 'sd798;
        'd355: dout <= -'sd777;
        'd356: dout <= 'sd912;
        'd357: dout <= -'sd298;
        'd358: dout <= -'sd950;
        'd359: dout <= -'sd480;
        'd360: dout <= -'sd2257;
        'd361: dout <= 'sd1008;
        'd362: dout <= 'sd645;
        'd363: dout <= -'sd1670;
        'd364: dout <= 'sd2286;
        'd365: dout <= 'sd643;
        'd366: dout <= 'sd1635;
        'd367: dout <= 'sd2136;
        'd368: dout <= 'sd630;
        'd369: dout <= -'sd1424;
        'd370: dout <= -'sd1966;
        'd371: dout <= -'sd1829;
        'd372: dout <= -'sd258;
        'd373: dout <= -'sd2130;
        'd374: dout <= 'sd998;
        'd375: dout <= 'sd1537;
        'd376: dout <= -'sd1381;
        'd377: dout <= 'sd1075;
        'd378: dout <= -'sd430;
        'd379: dout <= 'sd958;
        'd380: dout <= 'sd2017;
        'd381: dout <= 'sd320;
        'd382: dout <= -'sd505;
        'd383: dout <= 'sd1806;
        'd384: dout <= -'sd1909;
        'd385: dout <= 'sd1742;
        'd386: dout <= 'sd1105;
        'd387: dout <= -'sd1158;
        'd388: dout <= -'sd842;
        'd389: dout <= 'sd2238;
        'd390: dout <= -'sd357;
        'd391: dout <= -'sd41;
        'd392: dout <= -'sd349;
        'd393: dout <= -'sd905;
        'd394: dout <= 'sd548;
        'd395: dout <= -'sd1032;
        'd396: dout <= -'sd894;
        'd397: dout <= 'sd3;
        'd398: dout <= 'sd322;
        'd399: dout <= -'sd2032;
        'd400: dout <= -'sd922;
        'd401: dout <= 'sd777;
        'd402: dout <= -'sd1995;
        'd403: dout <= -'sd1022;
        'd404: dout <= -'sd1720;
        'd405: dout <= 'sd2215;
        'd406: dout <= 'sd2004;
        'd407: dout <= 'sd2167;
        'd408: dout <= 'sd943;
        'd409: dout <= -'sd845;
        'd410: dout <= -'sd2137;
        'd411: dout <= -'sd530;
        'd412: dout <= -'sd963;
        'd413: dout <= 'sd1468;
        'd414: dout <= 'sd277;
        'd415: dout <= 'sd2140;
        'd416: dout <= -'sd1129;
        'd417: dout <= 'sd1747;
        'd418: dout <= -'sd2231;
        'd419: dout <= 'sd2166;
        'd420: dout <= -'sd523;
        'd421: dout <= 'sd1543;
        'd422: dout <= 'sd1483;
        'd423: dout <= -'sd1817;
        'd424: dout <= -'sd1229;
        'd425: dout <= 'sd320;
        'd426: dout <= -'sd1770;
        'd427: dout <= -'sd994;
        'd428: dout <= 'sd1844;
        'd429: dout <= -'sd1651;
        'd430: dout <= -'sd1386;
        'd431: dout <= -'sd1310;
        'd432: dout <= -'sd36;
        'd433: dout <= 'sd1152;
        'd434: dout <= -'sd1264;
        'd435: dout <= 'sd555;
        'd436: dout <= 'sd1508;
        'd437: dout <= -'sd86;
        'd438: dout <= 'sd1448;
        'd439: dout <= -'sd2037;
        'd440: dout <= 'sd1961;
        'd441: dout <= -'sd2011;
        'd442: dout <= 'sd1216;
        'd443: dout <= 'sd507;
        'd444: dout <= -'sd1520;
        'd445: dout <= -'sd938;
        'd446: dout <= -'sd1255;
        'd447: dout <= 'sd1060;
        'd448: dout <= 'sd574;
        'd449: dout <= 'sd2218;
        'd450: dout <= -'sd1524;
        'd451: dout <= -'sd881;
        'd452: dout <= -'sd580;
        'd453: dout <= -'sd1215;
        'd454: dout <= 'sd719;
        'd455: dout <= 'sd2060;
        'd456: dout <= -'sd2160;
        'd457: dout <= -'sd1422;
        'd458: dout <= -'sd2166;
        'd459: dout <= 'sd403;
        'd460: dout <= 'sd1734;
        'd461: dout <= -'sd324;
        'd462: dout <= 'sd1203;
        'd463: dout <= 'sd263;
        'd464: dout <= -'sd2201;
        'd465: dout <= 'sd2188;
        'd466: dout <= 'sd1061;
        'd467: dout <= 'sd1844;
        'd468: dout <= -'sd354;
        'd469: dout <= 'sd1259;
        'd470: dout <= 'sd1788;
        'd471: dout <= 'sd1531;
        'd472: dout <= -'sd1787;
        'd473: dout <= -'sd207;
        'd474: dout <= -'sd1751;
        'd475: dout <= 'sd2229;
        'd476: dout <= 'sd773;
        'd477: dout <= 'sd406;
        'd478: dout <= -'sd970;
        'd479: dout <= 'sd122;
        'd480: dout <= 'sd2288;
        'd481: dout <= 'sd2237;
        'd482: dout <= 'sd316;
        'd483: dout <= -'sd550;
        'd484: dout <= 'sd1816;
        'd485: dout <= 'sd1962;
        'd486: dout <= 'sd2169;
        'd487: dout <= -'sd554;
        'd488: dout <= -'sd1936;
        'd489: dout <= 'sd514;
        'd490: dout <= -'sd748;
        'd491: dout <= -'sd154;
        'd492: dout <= 'sd1793;
        'd493: dout <= -'sd1561;
        'd494: dout <= 'sd1618;
        'd495: dout <= -'sd1015;
        'd496: dout <= 'sd618;
        'd497: dout <= 'sd1722;
        'd498: dout <= 'sd373;
        'd499: dout <= 'sd2107;
        'd500: dout <= 'sd643;
        'd501: dout <= -'sd614;
        'd502: dout <= 'sd14;
        'd503: dout <= -'sd753;
        'd504: dout <= -'sd1650;
        'd505: dout <= 'sd33;
        'd506: dout <= -'sd656;
        'd507: dout <= -'sd1826;
        'd508: dout <= -'sd1438;
        'd509: dout <= -'sd1982;
        'd510: dout <= 'sd1888;
        'd511: dout <= 'sd1666;
        'd512: dout <= 'sd556;
        'd513: dout <= -'sd1888;
        'd514: dout <= -'sd1850;
        'd515: dout <= 'sd1323;
        'd516: dout <= -'sd1146;
        'd517: dout <= 'sd267;
        'd518: dout <= 'sd160;
        'd519: dout <= -'sd1666;
        'd520: dout <= 'sd2237;
        'd521: dout <= -'sd1500;
        'd522: dout <= 'sd265;
        'd523: dout <= 'sd984;
        'd524: dout <= -'sd51;
        'd525: dout <= -'sd1973;
        'd526: dout <= 'sd478;
        'd527: dout <= -'sd76;
        'd528: dout <= 'sd67;
        'd529: dout <= 'sd807;
        'd530: dout <= -'sd1764;
        'd531: dout <= 'sd172;
        'd532: dout <= 'sd648;
        'd533: dout <= -'sd1851;
        'd534: dout <= -'sd813;
        'd535: dout <= -'sd734;
        'd536: dout <= 'sd609;
        'd537: dout <= -'sd87;
        'd538: dout <= 'sd1076;
        'd539: dout <= 'sd883;
        'd540: dout <= -'sd2107;
        'd541: dout <= -'sd534;
        'd542: dout <= -'sd1050;
        'd543: dout <= -'sd2112;
        'd544: dout <= 'sd661;
        'd545: dout <= -'sd76;
        'd546: dout <= 'sd1096;
        'd547: dout <= -'sd1252;
        'd548: dout <= -'sd1785;
        'd549: dout <= 'sd75;
        'd550: dout <= -'sd677;
        'd551: dout <= -'sd1039;
        'd552: dout <= -'sd430;
        'd553: dout <= 'sd1530;
        'd554: dout <= 'sd198;
        'd555: dout <= -'sd1300;
        'd556: dout <= 'sd1822;
        'd557: dout <= -'sd1703;
        'd558: dout <= 'sd34;
        'd559: dout <= 'sd317;
        'd560: dout <= 'sd1872;
        'd561: dout <= -'sd283;
        'd562: dout <= 'sd968;
        'd563: dout <= -'sd1526;
        'd564: dout <= -'sd195;
        'd565: dout <= -'sd2080;
        'd566: dout <= -'sd548;
        'd567: dout <= 'sd1511;
        'd568: dout <= -'sd942;
        'd569: dout <= 'sd692;
        'd570: dout <= -'sd1403;
        'd571: dout <= -'sd482;
        'd572: dout <= -'sd2071;
        'd573: dout <= -'sd340;
        'd574: dout <= 'sd981;
        'd575: dout <= 'sd1324;
        'd576: dout <= 'sd526;
        'd577: dout <= -'sd945;
        'd578: dout <= -'sd1464;
        'd579: dout <= 'sd1762;
        'd580: dout <= 'sd466;
        'd581: dout <= 'sd1451;
        'd582: dout <= -'sd1427;
        'd583: dout <= -'sd1849;
        'd584: dout <= 'sd1489;
        'd585: dout <= -'sd647;
        'd586: dout <= 'sd106;
        'd587: dout <= -'sd1566;
        'd588: dout <= 'sd1311;
        'd589: dout <= 'sd531;
        'd590: dout <= 'sd1849;
        'd591: dout <= -'sd812;
        'd592: dout <= -'sd202;
        'd593: dout <= -'sd1317;
        'd594: dout <= 'sd374;
        'd595: dout <= -'sd17;
        'd596: dout <= -'sd1067;
        'd597: dout <= -'sd1478;
        'd598: dout <= -'sd500;
        'd599: dout <= 'sd524;
        'd600: dout <= -'sd1748;
        'd601: dout <= -'sd1841;
        'd602: dout <= -'sd537;
        'd603: dout <= -'sd1216;
        'd604: dout <= -'sd1425;
        'd605: dout <= -'sd1004;
        'd606: dout <= -'sd1166;
        'd607: dout <= 'sd1981;
        'd608: dout <= -'sd1468;
        'd609: dout <= 'sd1588;
        'd610: dout <= -'sd150;
        'd611: dout <= -'sd789;
        'd612: dout <= 'sd1616;
        'd613: dout <= -'sd2024;
        'd614: dout <= -'sd213;
        'd615: dout <= 'sd1828;
        'd616: dout <= 'sd1395;
        'd617: dout <= 'sd1580;
        'd618: dout <= -'sd830;
        'd619: dout <= 'sd577;
        'd620: dout <= 'sd1157;
        'd621: dout <= -'sd497;
        'd622: dout <= 'sd1551;
        'd623: dout <= 'sd1673;
        'd624: dout <= -'sd1198;
        'd625: dout <= -'sd1101;
        'd626: dout <= -'sd1582;
        'd627: dout <= 'sd2288;
        'd628: dout <= -'sd521;
        'd629: dout <= 'sd1587;
        'd630: dout <= -'sd1310;
        'd631: dout <= -'sd1810;
        'd632: dout <= -'sd887;
        'd633: dout <= 'sd420;
        'd634: dout <= 'sd1692;
        'd635: dout <= 'sd2201;
        'd636: dout <= -'sd181;
        'd637: dout <= -'sd59;
        'd638: dout <= 'sd1627;
        'd639: dout <= -'sd992;
        'd640: dout <= 'sd2157;
        'd641: dout <= -'sd978;
        'd642: dout <= 'sd2138;
        'd643: dout <= -'sd1991;
        'd644: dout <= -'sd851;
        'd645: dout <= -'sd1955;
        'd646: dout <= -'sd391;
        'd647: dout <= -'sd2047;
        'd648: dout <= 'sd505;
        'd649: dout <= 'sd2199;
        'd650: dout <= -'sd1493;
        'd651: dout <= -'sd1912;
        'd652: dout <= -'sd2041;
        'd653: dout <= -'sd1402;
        'd654: dout <= -'sd1710;
        'd655: dout <= -'sd1771;
        'd656: dout <= 'sd2200;
        'd657: dout <= 'sd91;
        'd658: dout <= -'sd2239;
        'd659: dout <= -'sd405;
        'd660: dout <= 'sd2249;
        'd661: dout <= -'sd662;
        'd662: dout <= -'sd1048;
        'd663: dout <= -'sd411;
        'd664: dout <= 'sd1698;
        'd665: dout <= -'sd1476;
        'd666: dout <= 'sd536;
        'd667: dout <= -'sd1355;
        'd668: dout <= -'sd965;
        'd669: dout <= 'sd60;
        'd670: dout <= 'sd2210;
        'd671: dout <= -'sd772;
        'd672: dout <= -'sd371;
        'd673: dout <= -'sd1195;
        'd674: dout <= 'sd1926;
        'd675: dout <= 'sd1698;
        'd676: dout <= 'sd1713;
        'd677: dout <= -'sd909;
        'd678: dout <= 'sd221;
        'd679: dout <= 'sd499;
        'd680: dout <= -'sd1403;
        'd681: dout <= 'sd2044;
        'd682: dout <= 'sd404;
        'd683: dout <= -'sd109;
        'd684: dout <= 'sd376;
        'd685: dout <= -'sd1347;
        'd686: dout <= 'sd1311;
        'd687: dout <= -'sd1699;
        'd688: dout <= -'sd415;
        'd689: dout <= -'sd1272;
        'd690: dout <= -'sd2019;
        'd691: dout <= -'sd1752;
        'd692: dout <= 'sd1361;
        'd693: dout <= -'sd801;
        'd694: dout <= 'sd394;
        'd695: dout <= 'sd601;
        'd696: dout <= -'sd1770;
        'd697: dout <= 'sd412;
        'd698: dout <= 'sd562;
        'd699: dout <= -'sd1176;
        'd700: dout <= 'sd2038;
        'd701: dout <= -'sd516;
        'd702: dout <= -'sd2028;
        'd703: dout <= 'sd817;
        'd704: dout <= -'sd1362;
        'd705: dout <= -'sd195;
        'd706: dout <= 'sd1279;
        'd707: dout <= -'sd1489;
        'd708: dout <= 'sd2249;
        'd709: dout <= 'sd286;
        'd710: dout <= 'sd1717;
        'd711: dout <= 'sd1296;
        'd712: dout <= -'sd922;
        'd713: dout <= 'sd1413;
        'd714: dout <= -'sd1647;
        'd715: dout <= -'sd1865;
        'd716: dout <= -'sd655;
        'd717: dout <= 'sd1765;
        'd718: dout <= -'sd777;
        'd719: dout <= -'sd1176;
        'd720: dout <= 'sd291;
        'd721: dout <= 'sd1017;
        'd722: dout <= 'sd1019;
        'd723: dout <= -'sd937;
        'd724: dout <= -'sd195;
        'd725: dout <= 'sd1441;
        'd726: dout <= 'sd2090;
        'd727: dout <= 'sd1750;
        'd728: dout <= 'sd741;
        'd729: dout <= 'sd1031;
        'd730: dout <= -'sd1894;
        'd731: dout <= 'sd883;
        'd732: dout <= 'sd2211;
        'd733: dout <= -'sd2066;
        'd734: dout <= -'sd1056;
        'd735: dout <= -'sd350;
        'd736: dout <= 'sd503;
        'd737: dout <= 'sd230;
        'd738: dout <= -'sd1597;
        'd739: dout <= -'sd1572;
        'd740: dout <= 'sd59;
        'd741: dout <= 'sd1741;
        'd742: dout <= 'sd1371;
        'd743: dout <= -'sd675;
        'd744: dout <= -'sd561;
        'd745: dout <= -'sd1022;
        'd746: dout <= -'sd1812;
        'd747: dout <= 'sd1840;
        'd748: dout <= -'sd1803;
        'd749: dout <= 'sd1419;
        'd750: dout <= -'sd996;
        'd751: dout <= 'sd560;
        'd752: dout <= 'sd2116;
        'd753: dout <= -'sd867;
        'd754: dout <= 'sd545;
        'd755: dout <= 'sd1721;
        'd756: dout <= 'sd86;
        'd757: dout <= -'sd1042;
        'd758: dout <= -'sd1723;
        'd759: dout <= 'sd2223;
        'd760: dout <= -'sd130;
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module h_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [13:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'd0: dout <= -'sd2205;
        'd1: dout <= -'sd556;
        'd2: dout <= 'sd1047;
        'd3: dout <= -'sd877;
        'd4: dout <= -'sd309;
        'd5: dout <= 'sd676;
        'd6: dout <= -'sd124;
        'd7: dout <= 'sd1143;
        'd8: dout <= -'sd984;
        'd9: dout <= 'sd439;
        'd10: dout <= 'sd999;
        'd11: dout <= -'sd238;
        'd12: dout <= -'sd1941;
        'd13: dout <= 'sd1556;
        'd14: dout <= 'sd1746;
        'd15: dout <= -'sd2;
        'd16: dout <= 'sd2133;
        'd17: dout <= -'sd1076;
        'd18: dout <= -'sd1664;
        'd19: dout <= -'sd1349;
        'd20: dout <= -'sd864;
        'd21: dout <= 'sd762;
        'd22: dout <= 'sd144;
        'd23: dout <= -'sd2162;
        'd24: dout <= 'sd1892;
        'd25: dout <= 'sd936;
        'd26: dout <= -'sd1228;
        'd27: dout <= -'sd219;
        'd28: dout <= -'sd2074;
        'd29: dout <= -'sd791;
        'd30: dout <= 'sd1810;
        'd31: dout <= -'sd1806;
        'd32: dout <= 'sd1855;
        'd33: dout <= 'sd236;
        'd34: dout <= 'sd1236;
        'd35: dout <= 'sd464;
        'd36: dout <= -'sd1336;
        'd37: dout <= 'sd814;
        'd38: dout <= 'sd1506;
        'd39: dout <= -'sd1358;
        'd40: dout <= -'sd413;
        'd41: dout <= 'sd1939;
        'd42: dout <= -'sd1575;
        'd43: dout <= -'sd707;
        'd44: dout <= 'sd1505;
        'd45: dout <= 'sd2121;
        'd46: dout <= 'sd2069;
        'd47: dout <= 'sd1001;
        'd48: dout <= -'sd1341;
        'd49: dout <= -'sd86;
        'd50: dout <= -'sd2196;
        'd51: dout <= -'sd113;
        'd52: dout <= 'sd408;
        'd53: dout <= 'sd2050;
        'd54: dout <= -'sd1805;
        'd55: dout <= 'sd617;
        'd56: dout <= -'sd1717;
        'd57: dout <= 'sd336;
        'd58: dout <= -'sd1976;
        'd59: dout <= -'sd743;
        'd60: dout <= 'sd247;
        'd61: dout <= 'sd1810;
        'd62: dout <= -'sd1432;
        'd63: dout <= -'sd1741;
        'd64: dout <= -'sd891;
        'd65: dout <= 'sd2279;
        'd66: dout <= 'sd709;
        'd67: dout <= -'sd2183;
        'd68: dout <= 'sd2149;
        'd69: dout <= 'sd2031;
        'd70: dout <= -'sd1178;
        'd71: dout <= 'sd1459;
        'd72: dout <= 'sd0;
        'd73: dout <= -'sd981;
        'd74: dout <= 'sd495;
        'd75: dout <= 'sd492;
        'd76: dout <= -'sd882;
        'd77: dout <= -'sd1440;
        'd78: dout <= 'sd1201;
        'd79: dout <= -'sd202;
        'd80: dout <= -'sd1554;
        'd81: dout <= -'sd806;
        'd82: dout <= -'sd1271;
        'd83: dout <= -'sd1305;
        'd84: dout <= 'sd236;
        'd85: dout <= -'sd428;
        'd86: dout <= -'sd839;
        'd87: dout <= 'sd1372;
        'd88: dout <= 'sd1546;
        'd89: dout <= 'sd471;
        'd90: dout <= -'sd162;
        'd91: dout <= 'sd559;
        'd92: dout <= 'sd1585;
        'd93: dout <= 'sd8;
        'd94: dout <= 'sd1921;
        'd95: dout <= -'sd1506;
        'd96: dout <= 'sd176;
        'd97: dout <= -'sd799;
        'd98: dout <= 'sd833;
        'd99: dout <= -'sd1200;
        'd100: dout <= 'sd24;
        'd101: dout <= 'sd2264;
        'd102: dout <= 'sd785;
        'd103: dout <= 'sd1126;
        'd104: dout <= 'sd2106;
        'd105: dout <= 'sd1582;
        'd106: dout <= 'sd159;
        'd107: dout <= -'sd90;
        'd108: dout <= -'sd1600;
        'd109: dout <= 'sd561;
        'd110: dout <= 'sd2162;
        'd111: dout <= -'sd982;
        'd112: dout <= -'sd715;
        'd113: dout <= 'sd1544;
        'd114: dout <= -'sd1159;
        'd115: dout <= -'sd1108;
        'd116: dout <= 'sd1868;
        'd117: dout <= 'sd229;
        'd118: dout <= -'sd129;
        'd119: dout <= -'sd741;
        'd120: dout <= -'sd317;
        'd121: dout <= 'sd243;
        'd122: dout <= -'sd1113;
        'd123: dout <= 'sd349;
        'd124: dout <= -'sd270;
        'd125: dout <= 'sd438;
        'd126: dout <= 'sd1800;
        'd127: dout <= 'sd1536;
        'd128: dout <= -'sd261;
        'd129: dout <= 'sd724;
        'd130: dout <= -'sd876;
        'd131: dout <= 'sd1712;
        'd132: dout <= -'sd2220;
        'd133: dout <= 'sd1777;
        'd134: dout <= -'sd1991;
        'd135: dout <= 'sd1048;
        'd136: dout <= -'sd905;
        'd137: dout <= -'sd2093;
        'd138: dout <= -'sd1107;
        'd139: dout <= 'sd77;
        'd140: dout <= -'sd1614;
        'd141: dout <= 'sd1576;
        'd142: dout <= -'sd1762;
        'd143: dout <= -'sd330;
        'd144: dout <= -'sd819;
        'd145: dout <= -'sd1790;
        'd146: dout <= -'sd5;
        'd147: dout <= 'sd390;
        'd148: dout <= 'sd541;
        'd149: dout <= -'sd2268;
        'd150: dout <= -'sd2253;
        'd151: dout <= -'sd355;
        'd152: dout <= -'sd1701;
        'd153: dout <= 'sd2192;
        'd154: dout <= 'sd508;
        'd155: dout <= -'sd1024;
        'd156: dout <= -'sd2253;
        'd157: dout <= -'sd2217;
        'd158: dout <= 'sd276;
        'd159: dout <= 'sd456;
        'd160: dout <= 'sd752;
        'd161: dout <= 'sd1783;
        'd162: dout <= 'sd167;
        'd163: dout <= -'sd1900;
        'd164: dout <= 'sd1556;
        'd165: dout <= 'sd81;
        'd166: dout <= -'sd508;
        'd167: dout <= -'sd1511;
        'd168: dout <= -'sd2133;
        'd169: dout <= -'sd1744;
        'd170: dout <= 'sd1391;
        'd171: dout <= 'sd1313;
        'd172: dout <= -'sd2284;
        'd173: dout <= -'sd363;
        'd174: dout <= 'sd762;
        'd175: dout <= 'sd665;
        'd176: dout <= -'sd191;
        'd177: dout <= -'sd990;
        'd178: dout <= 'sd742;
        'd179: dout <= 'sd1354;
        'd180: dout <= 'sd914;
        'd181: dout <= -'sd1662;
        'd182: dout <= -'sd1654;
        'd183: dout <= 'sd1029;
        'd184: dout <= -'sd478;
        'd185: dout <= -'sd927;
        'd186: dout <= -'sd1832;
        'd187: dout <= 'sd1254;
        'd188: dout <= 'sd1582;
        'd189: dout <= 'sd519;
        'd190: dout <= 'sd1986;
        'd191: dout <= 'sd1756;
        'd192: dout <= 'sd2157;
        'd193: dout <= -'sd2267;
        'd194: dout <= 'sd1190;
        'd195: dout <= 'sd1440;
        'd196: dout <= -'sd2202;
        'd197: dout <= 'sd631;
        'd198: dout <= -'sd896;
        'd199: dout <= 'sd1123;
        'd200: dout <= -'sd1224;
        'd201: dout <= 'sd1244;
        'd202: dout <= 'sd1054;
        'd203: dout <= -'sd2032;
        'd204: dout <= 'sd1810;
        'd205: dout <= -'sd1107;
        'd206: dout <= 'sd132;
        'd207: dout <= 'sd1256;
        'd208: dout <= -'sd576;
        'd209: dout <= -'sd170;
        'd210: dout <= -'sd1003;
        'd211: dout <= -'sd1220;
        'd212: dout <= 'sd919;
        'd213: dout <= -'sd571;
        'd214: dout <= -'sd428;
        'd215: dout <= -'sd165;
        'd216: dout <= -'sd2221;
        'd217: dout <= -'sd521;
        'd218: dout <= 'sd2046;
        'd219: dout <= -'sd319;
        'd220: dout <= 'sd929;
        'd221: dout <= -'sd1015;
        'd222: dout <= 'sd1385;
        'd223: dout <= -'sd2062;
        'd224: dout <= -'sd786;
        'd225: dout <= 'sd835;
        'd226: dout <= 'sd1883;
        'd227: dout <= -'sd1576;
        'd228: dout <= 'sd165;
        'd229: dout <= -'sd1601;
        'd230: dout <= -'sd77;
        'd231: dout <= 'sd1432;
        'd232: dout <= 'sd1066;
        'd233: dout <= -'sd123;
        'd234: dout <= 'sd40;
        'd235: dout <= 'sd191;
        'd236: dout <= -'sd2084;
        'd237: dout <= 'sd551;
        'd238: dout <= 'sd2250;
        'd239: dout <= 'sd841;
        'd240: dout <= -'sd1008;
        'd241: dout <= 'sd1640;
        'd242: dout <= 'sd1323;
        'd243: dout <= 'sd2197;
        'd244: dout <= -'sd2131;
        'd245: dout <= 'sd2213;
        'd246: dout <= 'sd1742;
        'd247: dout <= -'sd2035;
        'd248: dout <= -'sd2004;
        'd249: dout <= 'sd45;
        'd250: dout <= -'sd354;
        'd251: dout <= 'sd477;
        'd252: dout <= -'sd1116;
        'd253: dout <= 'sd1142;
        'd254: dout <= -'sd462;
        'd255: dout <= 'sd1485;
        'd256: dout <= 'sd2222;
        'd257: dout <= -'sd751;
        'd258: dout <= 'sd177;
        'd259: dout <= 'sd2179;
        'd260: dout <= -'sd2036;
        'd261: dout <= 'sd82;
        'd262: dout <= -'sd1679;
        'd263: dout <= 'sd2072;
        'd264: dout <= 'sd498;
        'd265: dout <= -'sd1684;
        'd266: dout <= 'sd2198;
        'd267: dout <= 'sd1781;
        'd268: dout <= 'sd709;
        'd269: dout <= 'sd1822;
        'd270: dout <= 'sd2179;
        'd271: dout <= -'sd355;
        'd272: dout <= 'sd836;
        'd273: dout <= -'sd1297;
        'd274: dout <= -'sd112;
        'd275: dout <= 'sd566;
        'd276: dout <= 'sd1866;
        'd277: dout <= 'sd957;
        'd278: dout <= 'sd294;
        'd279: dout <= 'sd2173;
        'd280: dout <= -'sd1286;
        'd281: dout <= 'sd417;
        'd282: dout <= -'sd463;
        'd283: dout <= -'sd1401;
        'd284: dout <= -'sd739;
        'd285: dout <= -'sd1066;
        'd286: dout <= -'sd674;
        'd287: dout <= -'sd1771;
        'd288: dout <= 'sd1968;
        'd289: dout <= 'sd574;
        'd290: dout <= 'sd581;
        'd291: dout <= 'sd1060;
        'd292: dout <= 'sd878;
        'd293: dout <= -'sd631;
        'd294: dout <= 'sd116;
        'd295: dout <= 'sd181;
        'd296: dout <= -'sd871;
        'd297: dout <= 'sd1512;
        'd298: dout <= 'sd1153;
        'd299: dout <= -'sd932;
        'd300: dout <= -'sd966;
        'd301: dout <= 'sd2038;
        'd302: dout <= 'sd699;
        'd303: dout <= 'sd1199;
        'd304: dout <= 'sd2152;
        'd305: dout <= -'sd1798;
        'd306: dout <= 'sd1585;
        'd307: dout <= -'sd899;
        'd308: dout <= -'sd915;
        'd309: dout <= -'sd1064;
        'd310: dout <= 'sd1798;
        'd311: dout <= 'sd520;
        'd312: dout <= -'sd261;
        'd313: dout <= 'sd305;
        'd314: dout <= 'sd798;
        'd315: dout <= 'sd1542;
        'd316: dout <= 'sd2090;
        'd317: dout <= -'sd1086;
        'd318: dout <= -'sd1920;
        'd319: dout <= 'sd1782;
        'd320: dout <= 'sd1139;
        'd321: dout <= 'sd2222;
        'd322: dout <= -'sd1045;
        'd323: dout <= -'sd389;
        'd324: dout <= 'sd256;
        'd325: dout <= 'sd721;
        'd326: dout <= -'sd277;
        'd327: dout <= -'sd1988;
        'd328: dout <= 'sd1566;
        'd329: dout <= -'sd1955;
        'd330: dout <= -'sd1858;
        'd331: dout <= 'sd82;
        'd332: dout <= -'sd1726;
        'd333: dout <= -'sd1794;
        'd334: dout <= -'sd1039;
        'd335: dout <= 'sd832;
        'd336: dout <= -'sd1918;
        'd337: dout <= 'sd1428;
        'd338: dout <= -'sd498;
        'd339: dout <= -'sd28;
        'd340: dout <= 'sd86;
        'd341: dout <= -'sd631;
        'd342: dout <= -'sd364;
        'd343: dout <= 'sd332;
        'd344: dout <= 'sd17;
        'd345: dout <= 'sd1305;
        'd346: dout <= 'sd495;
        'd347: dout <= 'sd1838;
        'd348: dout <= 'sd306;
        'd349: dout <= -'sd760;
        'd350: dout <= -'sd2277;
        'd351: dout <= -'sd2156;
        'd352: dout <= 'sd243;
        'd353: dout <= 'sd1605;
        'd354: dout <= -'sd975;
        'd355: dout <= -'sd114;
        'd356: dout <= 'sd237;
        'd357: dout <= 'sd69;
        'd358: dout <= 'sd1266;
        'd359: dout <= -'sd510;
        'd360: dout <= -'sd356;
        'd361: dout <= 'sd583;
        'd362: dout <= -'sd2222;
        'd363: dout <= -'sd2125;
        'd364: dout <= 'sd26;
        'd365: dout <= 'sd220;
        'd366: dout <= 'sd177;
        'd367: dout <= -'sd1090;
        'd368: dout <= -'sd1598;
        'd369: dout <= 'sd2080;
        'd370: dout <= 'sd1792;
        'd371: dout <= -'sd18;
        'd372: dout <= -'sd2259;
        'd373: dout <= 'sd1901;
        'd374: dout <= 'sd2033;
        'd375: dout <= -'sd598;
        'd376: dout <= 'sd1670;
        'd377: dout <= 'sd1792;
        'd378: dout <= 'sd2270;
        'd379: dout <= 'sd926;
        'd380: dout <= -'sd1951;
        'd381: dout <= -'sd1665;
        'd382: dout <= -'sd52;
        'd383: dout <= -'sd988;
        'd384: dout <= -'sd2221;
        'd385: dout <= -'sd2092;
        'd386: dout <= -'sd1743;
        'd387: dout <= -'sd1611;
        'd388: dout <= -'sd1797;
        'd389: dout <= -'sd1469;
        'd390: dout <= 'sd1294;
        'd391: dout <= 'sd1405;
        'd392: dout <= -'sd500;
        'd393: dout <= -'sd1239;
        'd394: dout <= -'sd1551;
        'd395: dout <= 'sd2147;
        'd396: dout <= 'sd1117;
        'd397: dout <= -'sd2088;
        'd398: dout <= -'sd1760;
        'd399: dout <= -'sd1483;
        'd400: dout <= 'sd1323;
        'd401: dout <= -'sd2225;
        'd402: dout <= 'sd759;
        'd403: dout <= -'sd384;
        'd404: dout <= 'sd1582;
        'd405: dout <= 'sd1655;
        'd406: dout <= -'sd305;
        'd407: dout <= 'sd104;
        'd408: dout <= 'sd2115;
        'd409: dout <= -'sd2282;
        'd410: dout <= -'sd1644;
        'd411: dout <= -'sd134;
        'd412: dout <= -'sd1420;
        'd413: dout <= -'sd2180;
        'd414: dout <= -'sd2134;
        'd415: dout <= -'sd549;
        'd416: dout <= -'sd1160;
        'd417: dout <= -'sd137;
        'd418: dout <= 'sd432;
        'd419: dout <= -'sd2028;
        'd420: dout <= 'sd905;
        'd421: dout <= -'sd1321;
        'd422: dout <= 'sd529;
        'd423: dout <= -'sd458;
        'd424: dout <= 'sd1097;
        'd425: dout <= -'sd450;
        'd426: dout <= -'sd1576;
        'd427: dout <= 'sd383;
        'd428: dout <= 'sd800;
        'd429: dout <= 'sd759;
        'd430: dout <= 'sd794;
        'd431: dout <= 'sd1008;
        'd432: dout <= 'sd1248;
        'd433: dout <= -'sd1976;
        'd434: dout <= 'sd197;
        'd435: dout <= -'sd1997;
        'd436: dout <= -'sd2118;
        'd437: dout <= -'sd1209;
        'd438: dout <= 'sd58;
        'd439: dout <= -'sd1929;
        'd440: dout <= -'sd1647;
        'd441: dout <= -'sd1002;
        'd442: dout <= -'sd811;
        'd443: dout <= 'sd1985;
        'd444: dout <= -'sd1613;
        'd445: dout <= 'sd1573;
        'd446: dout <= -'sd2215;
        'd447: dout <= 'sd936;
        'd448: dout <= 'sd2049;
        'd449: dout <= -'sd2096;
        'd450: dout <= 'sd750;
        'd451: dout <= 'sd602;
        'd452: dout <= -'sd1990;
        'd453: dout <= 'sd1368;
        'd454: dout <= 'sd2100;
        'd455: dout <= 'sd1284;
        'd456: dout <= 'sd980;
        'd457: dout <= 'sd1414;
        'd458: dout <= -'sd264;
        'd459: dout <= 'sd155;
        'd460: dout <= 'sd125;
        'd461: dout <= 'sd2110;
        'd462: dout <= -'sd1445;
        'd463: dout <= -'sd296;
        'd464: dout <= -'sd257;
        'd465: dout <= -'sd467;
        'd466: dout <= 'sd1793;
        'd467: dout <= -'sd1809;
        'd468: dout <= 'sd1764;
        'd469: dout <= 'sd1746;
        'd470: dout <= -'sd987;
        'd471: dout <= 'sd888;
        'd472: dout <= 'sd1837;
        'd473: dout <= -'sd1498;
        'd474: dout <= -'sd205;
        'd475: dout <= -'sd421;
        'd476: dout <= 'sd743;
        'd477: dout <= -'sd552;
        'd478: dout <= 'sd450;
        'd479: dout <= -'sd678;
        'd480: dout <= -'sd1697;
        'd481: dout <= -'sd1215;
        'd482: dout <= -'sd2007;
        'd483: dout <= 'sd2175;
        'd484: dout <= 'sd2244;
        'd485: dout <= -'sd718;
        'd486: dout <= 'sd801;
        'd487: dout <= 'sd2118;
        'd488: dout <= 'sd294;
        'd489: dout <= 'sd1901;
        'd490: dout <= 'sd455;
        'd491: dout <= -'sd1292;
        'd492: dout <= 'sd2231;
        'd493: dout <= -'sd578;
        'd494: dout <= 'sd1435;
        'd495: dout <= 'sd1294;
        'd496: dout <= 'sd1868;
        'd497: dout <= 'sd458;
        'd498: dout <= -'sd297;
        'd499: dout <= 'sd1941;
        'd500: dout <= 'sd589;
        'd501: dout <= 'sd69;
        'd502: dout <= -'sd1428;
        'd503: dout <= -'sd1293;
        'd504: dout <= -'sd947;
        'd505: dout <= 'sd647;
        'd506: dout <= 'sd17;
        'd507: dout <= -'sd594;
        'd508: dout <= 'sd703;
        'd509: dout <= 'sd1290;
        'd510: dout <= 'sd1154;
        'd511: dout <= -'sd1401;
        'd512: dout <= -'sd960;
        'd513: dout <= -'sd1386;
        'd514: dout <= -'sd1596;
        'd515: dout <= -'sd1788;
        'd516: dout <= 'sd15;
        'd517: dout <= -'sd157;
        'd518: dout <= 'sd626;
        'd519: dout <= 'sd833;
        'd520: dout <= -'sd2031;
        'd521: dout <= 'sd179;
        'd522: dout <= 'sd1773;
        'd523: dout <= -'sd2284;
        'd524: dout <= -'sd1195;
        'd525: dout <= -'sd1091;
        'd526: dout <= 'sd889;
        'd527: dout <= -'sd1913;
        'd528: dout <= 'sd372;
        'd529: dout <= 'sd774;
        'd530: dout <= 'sd1279;
        'd531: dout <= -'sd186;
        'd532: dout <= -'sd187;
        'd533: dout <= -'sd1149;
        'd534: dout <= 'sd1195;
        'd535: dout <= 'sd253;
        'd536: dout <= -'sd1263;
        'd537: dout <= 'sd1361;
        'd538: dout <= -'sd2182;
        'd539: dout <= -'sd90;
        'd540: dout <= 'sd73;
        'd541: dout <= -'sd923;
        'd542: dout <= 'sd448;
        'd543: dout <= 'sd634;
        'd544: dout <= -'sd2050;
        'd545: dout <= 'sd692;
        'd546: dout <= 'sd1162;
        'd547: dout <= -'sd2041;
        'd548: dout <= -'sd660;
        'd549: dout <= 'sd148;
        'd550: dout <= 'sd175;
        'd551: dout <= 'sd520;
        'd552: dout <= 'sd1800;
        'd553: dout <= -'sd864;
        'd554: dout <= 'sd695;
        'd555: dout <= 'sd1285;
        'd556: dout <= 'sd942;
        'd557: dout <= 'sd2264;
        'd558: dout <= -'sd107;
        'd559: dout <= 'sd954;
        'd560: dout <= -'sd775;
        'd561: dout <= 'sd1721;
        'd562: dout <= 'sd1276;
        'd563: dout <= -'sd969;
        'd564: dout <= -'sd698;
        'd565: dout <= -'sd1111;
        'd566: dout <= 'sd756;
        'd567: dout <= -'sd1392;
        'd568: dout <= -'sd561;
        'd569: dout <= 'sd1884;
        'd570: dout <= 'sd401;
        'd571: dout <= -'sd1827;
        'd572: dout <= 'sd45;
        'd573: dout <= -'sd894;
        'd574: dout <= -'sd1877;
        'd575: dout <= 'sd1140;
        'd576: dout <= 'sd574;
        'd577: dout <= 'sd1533;
        'd578: dout <= 'sd1552;
        'd579: dout <= 'sd411;
        'd580: dout <= 'sd2060;
        'd581: dout <= -'sd1764;
        'd582: dout <= -'sd1641;
        'd583: dout <= 'sd2151;
        'd584: dout <= 'sd499;
        'd585: dout <= 'sd1046;
        'd586: dout <= 'sd1016;
        'd587: dout <= -'sd966;
        'd588: dout <= -'sd2291;
        'd589: dout <= 'sd801;
        'd590: dout <= 'sd1688;
        'd591: dout <= -'sd389;
        'd592: dout <= 'sd325;
        'd593: dout <= -'sd1411;
        'd594: dout <= -'sd140;
        'd595: dout <= 'sd733;
        'd596: dout <= -'sd766;
        'd597: dout <= 'sd816;
        'd598: dout <= -'sd764;
        'd599: dout <= -'sd1057;
        'd600: dout <= 'sd2011;
        'd601: dout <= 'sd1066;
        'd602: dout <= -'sd499;
        'd603: dout <= 'sd700;
        'd604: dout <= 'sd1040;
        'd605: dout <= 'sd290;
        'd606: dout <= -'sd715;
        'd607: dout <= 'sd1641;
        'd608: dout <= 'sd632;
        'd609: dout <= 'sd2118;
        'd610: dout <= 'sd1156;
        'd611: dout <= 'sd1908;
        'd612: dout <= -'sd351;
        'd613: dout <= 'sd2015;
        'd614: dout <= -'sd2053;
        'd615: dout <= 'sd1362;
        'd616: dout <= -'sd1409;
        'd617: dout <= 'sd342;
        'd618: dout <= -'sd260;
        'd619: dout <= -'sd1502;
        'd620: dout <= 'sd1388;
        'd621: dout <= 'sd1001;
        'd622: dout <= 'sd1093;
        'd623: dout <= 'sd859;
        'd624: dout <= -'sd2199;
        'd625: dout <= -'sd1488;
        'd626: dout <= -'sd2070;
        'd627: dout <= 'sd1508;
        'd628: dout <= 'sd1802;
        'd629: dout <= 'sd1397;
        'd630: dout <= -'sd515;
        'd631: dout <= 'sd2182;
        'd632: dout <= -'sd411;
        'd633: dout <= 'sd946;
        'd634: dout <= -'sd1496;
        'd635: dout <= -'sd496;
        'd636: dout <= 'sd1397;
        'd637: dout <= -'sd320;
        'd638: dout <= 'sd183;
        'd639: dout <= 'sd870;
        'd640: dout <= 'sd748;
        'd641: dout <= -'sd2073;
        'd642: dout <= 'sd11;
        'd643: dout <= -'sd636;
        'd644: dout <= -'sd640;
        'd645: dout <= -'sd469;
        'd646: dout <= -'sd1629;
        'd647: dout <= -'sd1518;
        'd648: dout <= 'sd1840;
        'd649: dout <= -'sd1628;
        'd650: dout <= 'sd2068;
        'd651: dout <= 'sd134;
        'd652: dout <= -'sd2131;
        'd653: dout <= 'sd1940;
        'd654: dout <= 'sd709;
        'd655: dout <= 'sd1741;
        'd656: dout <= -'sd1058;
        'd657: dout <= 'sd1247;
        'd658: dout <= -'sd2282;
        'd659: dout <= -'sd1261;
        'd660: dout <= 'sd1433;
        'd661: dout <= 'sd242;
        'd662: dout <= 'sd844;
        'd663: dout <= 'sd2176;
        'd664: dout <= -'sd2269;
        'd665: dout <= 'sd473;
        'd666: dout <= 'sd999;
        'd667: dout <= 'sd2155;
        'd668: dout <= 'sd1186;
        'd669: dout <= 'sd632;
        'd670: dout <= 'sd1521;
        'd671: dout <= -'sd1041;
        'd672: dout <= 'sd313;
        'd673: dout <= -'sd1750;
        'd674: dout <= -'sd22;
        'd675: dout <= -'sd1488;
        'd676: dout <= -'sd1557;
        'd677: dout <= 'sd1298;
        'd678: dout <= 'sd1820;
        'd679: dout <= 'sd2139;
        'd680: dout <= 'sd739;
        'd681: dout <= -'sd592;
        'd682: dout <= -'sd816;
        'd683: dout <= 'sd377;
        'd684: dout <= -'sd1884;
        'd685: dout <= -'sd386;
        'd686: dout <= -'sd2269;
        'd687: dout <= 'sd1826;
        'd688: dout <= -'sd816;
        'd689: dout <= -'sd812;
        'd690: dout <= 'sd1777;
        'd691: dout <= 'sd1087;
        'd692: dout <= 'sd2277;
        'd693: dout <= 'sd1244;
        'd694: dout <= 'sd1301;
        'd695: dout <= 'sd1082;
        'd696: dout <= -'sd170;
        'd697: dout <= 'sd1628;
        'd698: dout <= 'sd1143;
        'd699: dout <= 'sd541;
        'd700: dout <= 'sd314;
        'd701: dout <= 'sd1263;
        'd702: dout <= 'sd1613;
        'd703: dout <= 'sd678;
        'd704: dout <= 'sd319;
        'd705: dout <= -'sd437;
        'd706: dout <= -'sd1696;
        'd707: dout <= 'sd1785;
        'd708: dout <= -'sd2078;
        'd709: dout <= -'sd100;
        'd710: dout <= -'sd1482;
        'd711: dout <= -'sd891;
        'd712: dout <= -'sd2295;
        'd713: dout <= -'sd1000;
        'd714: dout <= -'sd73;
        'd715: dout <= -'sd375;
        'd716: dout <= -'sd1271;
        'd717: dout <= 'sd685;
        'd718: dout <= 'sd1140;
        'd719: dout <= -'sd364;
        'd720: dout <= -'sd226;
        'd721: dout <= -'sd1441;
        'd722: dout <= 'sd526;
        'd723: dout <= -'sd2114;
        'd724: dout <= 'sd1822;
        'd725: dout <= -'sd1872;
        'd726: dout <= 'sd288;
        'd727: dout <= -'sd992;
        'd728: dout <= 'sd1665;
        'd729: dout <= 'sd570;
        'd730: dout <= 'sd407;
        'd731: dout <= -'sd544;
        'd732: dout <= -'sd465;
        'd733: dout <= -'sd20;
        'd734: dout <= -'sd1624;
        'd735: dout <= -'sd244;
        'd736: dout <= -'sd439;
        'd737: dout <= 'sd1654;
        'd738: dout <= 'sd1121;
        'd739: dout <= -'sd1797;
        'd740: dout <= 'sd2279;
        'd741: dout <= -'sd2076;
        'd742: dout <= 'sd1762;
        'd743: dout <= -'sd1717;
        'd744: dout <= 'sd999;
        'd745: dout <= -'sd674;
        'd746: dout <= -'sd489;
        'd747: dout <= -'sd1178;
        'd748: dout <= -'sd1492;
        'd749: dout <= -'sd972;
        'd750: dout <= -'sd418;
        'd751: dout <= -'sd1596;
        'd752: dout <= 'sd541;
        'd753: dout <= -'sd303;
        'd754: dout <= 'sd2134;
        'd755: dout <= -'sd1864;
        'd756: dout <= 'sd2185;
        'd757: dout <= 'sd1325;
        'd758: dout <= -'sd1353;
        'd759: dout <= 'sd1095;
        'd760: dout <= -'sd2242;
        'd761: dout <= -'sd1375;
        'd762: dout <= -'sd623;
        'd763: dout <= -'sd1999;
        'd764: dout <= -'sd526;
        'd765: dout <= -'sd1566;
        'd766: dout <= 'sd699;
        'd767: dout <= -'sd2040;
        'd768: dout <= -'sd1130;
        'd769: dout <= -'sd976;
        'd770: dout <= 'sd1787;
        'd771: dout <= -'sd959;
        'd772: dout <= -'sd111;
        'd773: dout <= -'sd2193;
        'd774: dout <= -'sd948;
        'd775: dout <= 'sd1500;
        'd776: dout <= -'sd1247;
        'd777: dout <= 'sd324;
        'd778: dout <= -'sd16;
        'd779: dout <= 'sd1546;
        'd780: dout <= 'sd1495;
        'd781: dout <= 'sd1050;
        'd782: dout <= 'sd1525;
        'd783: dout <= 'sd750;
        'd784: dout <= -'sd500;
        'd785: dout <= -'sd1779;
        'd786: dout <= -'sd701;
        'd787: dout <= -'sd1385;
        'd788: dout <= -'sd1302;
        'd789: dout <= 'sd1065;
        'd790: dout <= 'sd1731;
        'd791: dout <= -'sd605;
        'd792: dout <= -'sd736;
        'd793: dout <= -'sd1650;
        'd794: dout <= -'sd1205;
        'd795: dout <= 'sd2179;
        'd796: dout <= -'sd2198;
        'd797: dout <= 'sd1588;
        'd798: dout <= 'sd14;
        'd799: dout <= 'sd1431;
        'd800: dout <= 'sd367;
        'd801: dout <= -'sd97;
        'd802: dout <= -'sd1543;
        'd803: dout <= 'sd1548;
        'd804: dout <= -'sd917;
        'd805: dout <= 'sd1039;
        'd806: dout <= -'sd865;
        'd807: dout <= 'sd2233;
        'd808: dout <= 'sd808;
        'd809: dout <= -'sd1042;
        'd810: dout <= 'sd1635;
        'd811: dout <= -'sd578;
        'd812: dout <= 'sd1679;
        'd813: dout <= -'sd9;
        'd814: dout <= 'sd1366;
        'd815: dout <= -'sd1047;
        'd816: dout <= 'sd1713;
        'd817: dout <= -'sd2255;
        'd818: dout <= 'sd931;
        'd819: dout <= 'sd1905;
        'd820: dout <= 'sd2204;
        'd821: dout <= -'sd614;
        'd822: dout <= 'sd376;
        'd823: dout <= 'sd1009;
        'd824: dout <= 'sd745;
        'd825: dout <= -'sd1547;
        'd826: dout <= 'sd1294;
        'd827: dout <= -'sd494;
        'd828: dout <= -'sd1907;
        'd829: dout <= 'sd716;
        'd830: dout <= -'sd993;
        'd831: dout <= 'sd683;
        'd832: dout <= -'sd620;
        'd833: dout <= 'sd377;
        'd834: dout <= -'sd1940;
        'd835: dout <= -'sd2210;
        'd836: dout <= -'sd255;
        'd837: dout <= 'sd1283;
        'd838: dout <= -'sd100;
        'd839: dout <= 'sd1252;
        'd840: dout <= 'sd882;
        'd841: dout <= 'sd1513;
        'd842: dout <= 'sd1552;
        'd843: dout <= -'sd1260;
        'd844: dout <= 'sd77;
        'd845: dout <= -'sd1073;
        'd846: dout <= 'sd1153;
        'd847: dout <= -'sd1498;
        'd848: dout <= 'sd679;
        'd849: dout <= 'sd1480;
        'd850: dout <= -'sd1113;
        'd851: dout <= 'sd1221;
        'd852: dout <= 'sd947;
        'd853: dout <= 'sd1825;
        'd854: dout <= -'sd1534;
        'd855: dout <= -'sd2171;
        'd856: dout <= 'sd2060;
        'd857: dout <= -'sd1902;
        'd858: dout <= -'sd1002;
        'd859: dout <= -'sd914;
        'd860: dout <= -'sd367;
        'd861: dout <= -'sd263;
        'd862: dout <= 'sd1203;
        'd863: dout <= 'sd2014;
        'd864: dout <= -'sd608;
        'd865: dout <= 'sd986;
        'd866: dout <= 'sd45;
        'd867: dout <= 'sd604;
        'd868: dout <= -'sd1671;
        'd869: dout <= -'sd1092;
        'd870: dout <= 'sd588;
        'd871: dout <= -'sd1185;
        'd872: dout <= 'sd1782;
        'd873: dout <= 'sd1922;
        'd874: dout <= -'sd1343;
        'd875: dout <= -'sd719;
        'd876: dout <= 'sd323;
        'd877: dout <= 'sd2277;
        'd878: dout <= -'sd1525;
        'd879: dout <= -'sd443;
        'd880: dout <= 'sd608;
        'd881: dout <= 'sd702;
        'd882: dout <= 'sd95;
        'd883: dout <= 'sd578;
        'd884: dout <= 'sd484;
        'd885: dout <= 'sd2107;
        'd886: dout <= -'sd43;
        'd887: dout <= -'sd1471;
        'd888: dout <= -'sd1511;
        'd889: dout <= -'sd805;
        'd890: dout <= 'sd1270;
        'd891: dout <= 'sd819;
        'd892: dout <= -'sd2278;
        'd893: dout <= 'sd1414;
        'd894: dout <= 'sd851;
        'd895: dout <= -'sd46;
        'd896: dout <= 'sd110;
        'd897: dout <= -'sd188;
        'd898: dout <= -'sd1299;
        'd899: dout <= 'sd1806;
        'd900: dout <= -'sd727;
        'd901: dout <= 'sd152;
        'd902: dout <= -'sd28;
        'd903: dout <= -'sd1151;
        'd904: dout <= -'sd758;
        'd905: dout <= -'sd138;
        'd906: dout <= 'sd1887;
        'd907: dout <= -'sd100;
        'd908: dout <= -'sd2038;
        'd909: dout <= -'sd1872;
        'd910: dout <= -'sd2079;
        'd911: dout <= -'sd1319;
        'd912: dout <= 'sd482;
        'd913: dout <= -'sd1565;
        'd914: dout <= -'sd267;
        'd915: dout <= 'sd602;
        'd916: dout <= -'sd163;
        'd917: dout <= -'sd671;
        'd918: dout <= 'sd652;
        'd919: dout <= -'sd159;
        'd920: dout <= 'sd1950;
        'd921: dout <= 'sd845;
        'd922: dout <= 'sd478;
        'd923: dout <= 'sd828;
        'd924: dout <= -'sd1408;
        'd925: dout <= -'sd2177;
        'd926: dout <= -'sd973;
        'd927: dout <= 'sd518;
        'd928: dout <= 'sd1059;
        'd929: dout <= 'sd921;
        'd930: dout <= 'sd1942;
        'd931: dout <= 'sd1340;
        'd932: dout <= -'sd2144;
        'd933: dout <= 'sd141;
        'd934: dout <= -'sd1144;
        'd935: dout <= 'sd1934;
        'd936: dout <= -'sd748;
        'd937: dout <= 'sd85;
        'd938: dout <= 'sd1204;
        'd939: dout <= 'sd1157;
        'd940: dout <= -'sd2211;
        'd941: dout <= 'sd105;
        'd942: dout <= -'sd1898;
        'd943: dout <= -'sd1698;
        'd944: dout <= 'sd1072;
        'd945: dout <= -'sd2138;
        'd946: dout <= -'sd376;
        'd947: dout <= -'sd168;
        'd948: dout <= -'sd2221;
        'd949: dout <= 'sd2107;
        'd950: dout <= -'sd2290;
        'd951: dout <= -'sd2044;
        'd952: dout <= -'sd834;
        'd953: dout <= -'sd1597;
        'd954: dout <= 'sd442;
        'd955: dout <= -'sd1099;
        'd956: dout <= 'sd57;
        'd957: dout <= 'sd582;
        'd958: dout <= -'sd517;
        'd959: dout <= 'sd1759;
        'd960: dout <= -'sd1067;
        'd961: dout <= -'sd1273;
        'd962: dout <= 'sd1187;
        'd963: dout <= -'sd455;
        'd964: dout <= -'sd2209;
        'd965: dout <= 'sd200;
        'd966: dout <= 'sd2176;
        'd967: dout <= 'sd747;
        'd968: dout <= 'sd1730;
        'd969: dout <= -'sd232;
        'd970: dout <= 'sd815;
        'd971: dout <= -'sd49;
        'd972: dout <= -'sd1575;
        'd973: dout <= -'sd1284;
        'd974: dout <= 'sd1905;
        'd975: dout <= 'sd670;
        'd976: dout <= 'sd700;
        'd977: dout <= -'sd827;
        'd978: dout <= -'sd961;
        'd979: dout <= 'sd1124;
        'd980: dout <= 'sd80;
        'd981: dout <= 'sd1866;
        'd982: dout <= 'sd205;
        'd983: dout <= -'sd1598;
        'd984: dout <= 'sd2056;
        'd985: dout <= 'sd315;
        'd986: dout <= -'sd1338;
        'd987: dout <= 'sd1245;
        'd988: dout <= -'sd326;
        'd989: dout <= 'sd1125;
        'd990: dout <= 'sd1176;
        'd991: dout <= -'sd723;
        'd992: dout <= -'sd1761;
        'd993: dout <= -'sd1958;
        'd994: dout <= 'sd2026;
        'd995: dout <= 'sd1934;
        'd996: dout <= 'sd1169;
        'd997: dout <= 'sd1512;
        'd998: dout <= -'sd1604;
        'd999: dout <= 'sd778;
        'd1000: dout <= 'sd1681;
        'd1001: dout <= -'sd1193;
        'd1002: dout <= 'sd1361;
        'd1003: dout <= 'sd854;
        'd1004: dout <= 'sd177;
        'd1005: dout <= -'sd430;
        'd1006: dout <= -'sd701;
        'd1007: dout <= 'sd1420;
        'd1008: dout <= -'sd74;
        'd1009: dout <= -'sd1142;
        'd1010: dout <= -'sd1566;
        'd1011: dout <= -'sd1782;
        'd1012: dout <= -'sd2187;
        'd1013: dout <= -'sd1646;
        'd1014: dout <= -'sd1067;
        'd1015: dout <= -'sd1940;
        'd1016: dout <= -'sd2022;
        'd1017: dout <= -'sd207;
        'd1018: dout <= 'sd1440;
        'd1019: dout <= -'sd1630;
        'd1020: dout <= -'sd1914;
        'd1021: dout <= 'sd1774;
        'd1022: dout <= -'sd818;
        'd1023: dout <= 'sd1133;
        'd1024: dout <= 'sd143;
        'd1025: dout <= 'sd56;
        'd1026: dout <= -'sd1207;
        'd1027: dout <= 'sd1029;
        'd1028: dout <= -'sd916;
        'd1029: dout <= 'sd2123;
        'd1030: dout <= 'sd640;
        'd1031: dout <= -'sd1859;
        'd1032: dout <= -'sd230;
        'd1033: dout <= 'sd2060;
        'd1034: dout <= -'sd1101;
        'd1035: dout <= 'sd983;
        'd1036: dout <= 'sd1123;
        'd1037: dout <= -'sd347;
        'd1038: dout <= -'sd2051;
        'd1039: dout <= -'sd1764;
        'd1040: dout <= -'sd118;
        'd1041: dout <= 'sd1273;
        'd1042: dout <= -'sd1462;
        'd1043: dout <= 'sd1279;
        'd1044: dout <= 'sd2240;
        'd1045: dout <= -'sd142;
        'd1046: dout <= 'sd621;
        'd1047: dout <= -'sd1478;
        'd1048: dout <= 'sd480;
        'd1049: dout <= 'sd2149;
        'd1050: dout <= 'sd348;
        'd1051: dout <= -'sd700;
        'd1052: dout <= -'sd1619;
        'd1053: dout <= -'sd348;
        'd1054: dout <= -'sd1232;
        'd1055: dout <= -'sd101;
        'd1056: dout <= 'sd1081;
        'd1057: dout <= -'sd706;
        'd1058: dout <= 'sd380;
        'd1059: dout <= 'sd2140;
        'd1060: dout <= 'sd772;
        'd1061: dout <= -'sd2059;
        'd1062: dout <= 'sd804;
        'd1063: dout <= 'sd1392;
        'd1064: dout <= 'sd1288;
        'd1065: dout <= -'sd1117;
        'd1066: dout <= 'sd1774;
        'd1067: dout <= 'sd2169;
        'd1068: dout <= 'sd868;
        'd1069: dout <= 'sd1651;
        'd1070: dout <= 'sd1414;
        'd1071: dout <= -'sd1657;
        'd1072: dout <= 'sd2172;
        'd1073: dout <= 'sd567;
        'd1074: dout <= -'sd2289;
        'd1075: dout <= 'sd284;
        'd1076: dout <= 'sd1380;
        'd1077: dout <= -'sd348;
        'd1078: dout <= -'sd138;
        'd1079: dout <= 'sd142;
        'd1080: dout <= 'sd2214;
        'd1081: dout <= -'sd1157;
        'd1082: dout <= 'sd385;
        'd1083: dout <= 'sd154;
        'd1084: dout <= -'sd2148;
        'd1085: dout <= 'sd1163;
        'd1086: dout <= -'sd293;
        'd1087: dout <= -'sd193;
        'd1088: dout <= 'sd655;
        'd1089: dout <= -'sd1600;
        'd1090: dout <= -'sd1906;
        'd1091: dout <= -'sd61;
        'd1092: dout <= -'sd1133;
        'd1093: dout <= 'sd2204;
        'd1094: dout <= 'sd326;
        'd1095: dout <= -'sd510;
        'd1096: dout <= -'sd2151;
        'd1097: dout <= 'sd1942;
        'd1098: dout <= 'sd1597;
        'd1099: dout <= -'sd1279;
        'd1100: dout <= 'sd1032;
        'd1101: dout <= -'sd31;
        'd1102: dout <= 'sd101;
        'd1103: dout <= -'sd457;
        'd1104: dout <= -'sd628;
        'd1105: dout <= 'sd1843;
        'd1106: dout <= -'sd1352;
        'd1107: dout <= -'sd248;
        'd1108: dout <= 'sd41;
        'd1109: dout <= -'sd1227;
        'd1110: dout <= -'sd1370;
        'd1111: dout <= -'sd330;
        'd1112: dout <= -'sd546;
        'd1113: dout <= 'sd1565;
        'd1114: dout <= -'sd1581;
        'd1115: dout <= -'sd2178;
        'd1116: dout <= -'sd754;
        'd1117: dout <= 'sd217;
        'd1118: dout <= -'sd959;
        'd1119: dout <= 'sd1647;
        'd1120: dout <= -'sd1742;
        'd1121: dout <= 'sd1914;
        'd1122: dout <= 'sd163;
        'd1123: dout <= 'sd378;
        'd1124: dout <= -'sd1028;
        'd1125: dout <= 'sd62;
        'd1126: dout <= -'sd1724;
        'd1127: dout <= -'sd1908;
        'd1128: dout <= 'sd785;
        'd1129: dout <= -'sd1094;
        'd1130: dout <= -'sd1916;
        'd1131: dout <= -'sd1368;
        'd1132: dout <= -'sd1576;
        'd1133: dout <= -'sd2045;
        'd1134: dout <= 'sd1099;
        'd1135: dout <= 'sd656;
        'd1136: dout <= -'sd1430;
        'd1137: dout <= -'sd736;
        'd1138: dout <= 'sd1849;
        'd1139: dout <= 'sd1275;
        'd1140: dout <= 'sd1188;
        'd1141: dout <= -'sd1350;
        'd1142: dout <= -'sd1401;
        'd1143: dout <= -'sd2046;
        'd1144: dout <= 'sd1685;
        'd1145: dout <= 'sd2256;
        'd1146: dout <= -'sd1966;
        'd1147: dout <= 'sd1572;
        'd1148: dout <= -'sd1439;
        'd1149: dout <= 'sd1989;
        'd1150: dout <= -'sd1393;
        'd1151: dout <= 'sd1780;
        'd1152: dout <= 'sd2082;
        'd1153: dout <= 'sd227;
        'd1154: dout <= -'sd365;
        'd1155: dout <= 'sd924;
        'd1156: dout <= 'sd1422;
        'd1157: dout <= 'sd375;
        'd1158: dout <= 'sd847;
        'd1159: dout <= 'sd995;
        'd1160: dout <= 'sd1012;
        'd1161: dout <= -'sd1169;
        'd1162: dout <= -'sd1811;
        'd1163: dout <= -'sd1104;
        'd1164: dout <= -'sd187;
        'd1165: dout <= -'sd1083;
        'd1166: dout <= 'sd1182;
        'd1167: dout <= 'sd904;
        'd1168: dout <= 'sd1011;
        'd1169: dout <= -'sd1077;
        'd1170: dout <= 'sd1167;
        'd1171: dout <= -'sd80;
        'd1172: dout <= 'sd773;
        'd1173: dout <= 'sd892;
        'd1174: dout <= 'sd147;
        'd1175: dout <= 'sd1666;
        'd1176: dout <= -'sd315;
        'd1177: dout <= -'sd642;
        'd1178: dout <= -'sd1190;
        'd1179: dout <= 'sd1834;
        'd1180: dout <= 'sd1731;
        'd1181: dout <= -'sd2146;
        'd1182: dout <= -'sd265;
        'd1183: dout <= 'sd772;
        'd1184: dout <= 'sd2079;
        'd1185: dout <= 'sd1931;
        'd1186: dout <= -'sd562;
        'd1187: dout <= 'sd1287;
        'd1188: dout <= -'sd323;
        'd1189: dout <= 'sd1045;
        'd1190: dout <= 'sd242;
        'd1191: dout <= 'sd2205;
        'd1192: dout <= 'sd1049;
        'd1193: dout <= -'sd1791;
        'd1194: dout <= 'sd281;
        'd1195: dout <= -'sd218;
        'd1196: dout <= -'sd1945;
        'd1197: dout <= -'sd1278;
        'd1198: dout <= -'sd2267;
        'd1199: dout <= 'sd571;
        'd1200: dout <= 'sd22;
        'd1201: dout <= -'sd1647;
        'd1202: dout <= 'sd1058;
        'd1203: dout <= 'sd1991;
        'd1204: dout <= 'sd283;
        'd1205: dout <= -'sd647;
        'd1206: dout <= 'sd1778;
        'd1207: dout <= 'sd2241;
        'd1208: dout <= -'sd532;
        'd1209: dout <= 'sd602;
        'd1210: dout <= -'sd520;
        'd1211: dout <= 'sd1265;
        'd1212: dout <= -'sd1419;
        'd1213: dout <= 'sd1751;
        'd1214: dout <= -'sd2130;
        'd1215: dout <= 'sd730;
        'd1216: dout <= 'sd2256;
        'd1217: dout <= 'sd1346;
        'd1218: dout <= 'sd1711;
        'd1219: dout <= -'sd950;
        'd1220: dout <= 'sd489;
        'd1221: dout <= -'sd1710;
        'd1222: dout <= -'sd129;
        'd1223: dout <= 'sd1219;
        'd1224: dout <= 'sd1996;
        'd1225: dout <= -'sd402;
        'd1226: dout <= -'sd1182;
        'd1227: dout <= -'sd1435;
        'd1228: dout <= 'sd168;
        'd1229: dout <= 'sd2177;
        'd1230: dout <= 'sd1180;
        'd1231: dout <= -'sd770;
        'd1232: dout <= -'sd136;
        'd1233: dout <= 'sd108;
        'd1234: dout <= -'sd978;
        'd1235: dout <= -'sd637;
        'd1236: dout <= -'sd1706;
        'd1237: dout <= 'sd837;
        'd1238: dout <= 'sd687;
        'd1239: dout <= 'sd1405;
        'd1240: dout <= -'sd381;
        'd1241: dout <= -'sd1280;
        'd1242: dout <= 'sd1754;
        'd1243: dout <= 'sd2067;
        'd1244: dout <= 'sd969;
        'd1245: dout <= -'sd60;
        'd1246: dout <= 'sd988;
        'd1247: dout <= -'sd939;
        'd1248: dout <= 'sd1638;
        'd1249: dout <= -'sd966;
        'd1250: dout <= 'sd1217;
        'd1251: dout <= 'sd523;
        'd1252: dout <= -'sd869;
        'd1253: dout <= 'sd725;
        'd1254: dout <= -'sd712;
        'd1255: dout <= -'sd1925;
        'd1256: dout <= 'sd2090;
        'd1257: dout <= -'sd1190;
        'd1258: dout <= 'sd1433;
        'd1259: dout <= 'sd1178;
        'd1260: dout <= -'sd1082;
        'd1261: dout <= 'sd1640;
        'd1262: dout <= 'sd2193;
        'd1263: dout <= -'sd159;
        'd1264: dout <= -'sd765;
        'd1265: dout <= 'sd564;
        'd1266: dout <= -'sd1804;
        'd1267: dout <= -'sd917;
        'd1268: dout <= -'sd1099;
        'd1269: dout <= -'sd247;
        'd1270: dout <= 'sd1116;
        'd1271: dout <= -'sd399;
        'd1272: dout <= 'sd70;
        'd1273: dout <= -'sd201;
        'd1274: dout <= -'sd1459;
        'd1275: dout <= 'sd5;
        'd1276: dout <= 'sd528;
        'd1277: dout <= -'sd1123;
        'd1278: dout <= -'sd1875;
        'd1279: dout <= 'sd1792;
        'd1280: dout <= 'sd1715;
        'd1281: dout <= -'sd24;
        'd1282: dout <= 'sd399;
        'd1283: dout <= -'sd312;
        'd1284: dout <= 'sd649;
        'd1285: dout <= 'sd1558;
        'd1286: dout <= -'sd1015;
        'd1287: dout <= 'sd821;
        'd1288: dout <= 'sd201;
        'd1289: dout <= 'sd357;
        'd1290: dout <= 'sd118;
        'd1291: dout <= 'sd160;
        'd1292: dout <= -'sd78;
        'd1293: dout <= 'sd1985;
        'd1294: dout <= -'sd515;
        'd1295: dout <= 'sd900;
        'd1296: dout <= -'sd440;
        'd1297: dout <= 'sd1614;
        'd1298: dout <= 'sd985;
        'd1299: dout <= -'sd2071;
        'd1300: dout <= -'sd839;
        'd1301: dout <= 'sd900;
        'd1302: dout <= -'sd1660;
        'd1303: dout <= -'sd1608;
        'd1304: dout <= 'sd482;
        'd1305: dout <= 'sd639;
        'd1306: dout <= -'sd876;
        'd1307: dout <= -'sd702;
        'd1308: dout <= 'sd2160;
        'd1309: dout <= -'sd655;
        'd1310: dout <= -'sd836;
        'd1311: dout <= -'sd1131;
        'd1312: dout <= 'sd465;
        'd1313: dout <= -'sd953;
        'd1314: dout <= -'sd1085;
        'd1315: dout <= 'sd42;
        'd1316: dout <= 'sd109;
        'd1317: dout <= -'sd1806;
        'd1318: dout <= 'sd1078;
        'd1319: dout <= -'sd917;
        'd1320: dout <= -'sd1935;
        'd1321: dout <= 'sd1894;
        'd1322: dout <= -'sd45;
        'd1323: dout <= 'sd432;
        'd1324: dout <= 'sd958;
        'd1325: dout <= 'sd600;
        'd1326: dout <= -'sd1803;
        'd1327: dout <= -'sd1185;
        'd1328: dout <= -'sd518;
        'd1329: dout <= 'sd310;
        'd1330: dout <= 'sd986;
        'd1331: dout <= 'sd2205;
        'd1332: dout <= 'sd1434;
        'd1333: dout <= -'sd1815;
        'd1334: dout <= 'sd1972;
        'd1335: dout <= -'sd927;
        'd1336: dout <= -'sd778;
        'd1337: dout <= -'sd1001;
        'd1338: dout <= -'sd1171;
        'd1339: dout <= 'sd479;
        'd1340: dout <= -'sd55;
        'd1341: dout <= -'sd904;
        'd1342: dout <= -'sd583;
        'd1343: dout <= 'sd2122;
        'd1344: dout <= 'sd1548;
        'd1345: dout <= 'sd1215;
        'd1346: dout <= -'sd1664;
        'd1347: dout <= 'sd399;
        'd1348: dout <= 'sd117;
        'd1349: dout <= -'sd908;
        'd1350: dout <= -'sd316;
        'd1351: dout <= 'sd359;
        'd1352: dout <= -'sd1290;
        'd1353: dout <= -'sd1497;
        'd1354: dout <= -'sd1949;
        'd1355: dout <= 'sd800;
        'd1356: dout <= -'sd391;
        'd1357: dout <= 'sd403;
        'd1358: dout <= 'sd1419;
        'd1359: dout <= 'sd2039;
        'd1360: dout <= -'sd1290;
        'd1361: dout <= 'sd310;
        'd1362: dout <= 'sd2109;
        'd1363: dout <= -'sd1998;
        'd1364: dout <= -'sd916;
        'd1365: dout <= -'sd1075;
        'd1366: dout <= -'sd1328;
        'd1367: dout <= -'sd1503;
        'd1368: dout <= 'sd443;
        'd1369: dout <= -'sd1452;
        'd1370: dout <= 'sd1148;
        'd1371: dout <= -'sd653;
        'd1372: dout <= 'sd2288;
        'd1373: dout <= -'sd1586;
        'd1374: dout <= 'sd403;
        'd1375: dout <= 'sd2161;
        'd1376: dout <= -'sd1181;
        'd1377: dout <= 'sd1124;
        'd1378: dout <= 'sd2028;
        'd1379: dout <= -'sd1363;
        'd1380: dout <= -'sd476;
        'd1381: dout <= -'sd909;
        'd1382: dout <= -'sd1853;
        'd1383: dout <= -'sd714;
        'd1384: dout <= -'sd1320;
        'd1385: dout <= -'sd2259;
        'd1386: dout <= 'sd1001;
        'd1387: dout <= -'sd456;
        'd1388: dout <= -'sd1163;
        'd1389: dout <= 'sd2239;
        'd1390: dout <= 'sd1333;
        'd1391: dout <= 'sd1388;
        'd1392: dout <= -'sd985;
        'd1393: dout <= 'sd2064;
        'd1394: dout <= -'sd526;
        'd1395: dout <= 'sd2218;
        'd1396: dout <= -'sd1201;
        'd1397: dout <= 'sd1104;
        'd1398: dout <= -'sd421;
        'd1399: dout <= 'sd758;
        'd1400: dout <= -'sd1200;
        'd1401: dout <= 'sd940;
        'd1402: dout <= 'sd1395;
        'd1403: dout <= -'sd1694;
        'd1404: dout <= 'sd1097;
        'd1405: dout <= 'sd2192;
        'd1406: dout <= -'sd2059;
        'd1407: dout <= -'sd1172;
        'd1408: dout <= -'sd620;
        'd1409: dout <= -'sd424;
        'd1410: dout <= 'sd1168;
        'd1411: dout <= -'sd1850;
        'd1412: dout <= -'sd1919;
        'd1413: dout <= 'sd1116;
        'd1414: dout <= 'sd257;
        'd1415: dout <= 'sd1158;
        'd1416: dout <= 'sd1288;
        'd1417: dout <= -'sd686;
        'd1418: dout <= 'sd1967;
        'd1419: dout <= 'sd618;
        'd1420: dout <= 'sd1736;
        'd1421: dout <= 'sd1880;
        'd1422: dout <= 'sd919;
        'd1423: dout <= 'sd71;
        'd1424: dout <= -'sd95;
        'd1425: dout <= 'sd1956;
        'd1426: dout <= 'sd1743;
        'd1427: dout <= -'sd280;
        'd1428: dout <= -'sd598;
        'd1429: dout <= 'sd475;
        'd1430: dout <= -'sd297;
        'd1431: dout <= -'sd1872;
        'd1432: dout <= 'sd1587;
        'd1433: dout <= -'sd1277;
        'd1434: dout <= 'sd1627;
        'd1435: dout <= -'sd698;
        'd1436: dout <= 'sd24;
        'd1437: dout <= 'sd1957;
        'd1438: dout <= 'sd1015;
        'd1439: dout <= 'sd855;
        'd1440: dout <= -'sd1376;
        'd1441: dout <= 'sd1583;
        'd1442: dout <= 'sd1033;
        'd1443: dout <= 'sd1401;
        'd1444: dout <= -'sd111;
        'd1445: dout <= 'sd953;
        'd1446: dout <= -'sd540;
        'd1447: dout <= -'sd922;
        'd1448: dout <= -'sd19;
        'd1449: dout <= -'sd2198;
        'd1450: dout <= -'sd2182;
        'd1451: dout <= -'sd679;
        'd1452: dout <= -'sd2250;
        'd1453: dout <= 'sd913;
        'd1454: dout <= -'sd110;
        'd1455: dout <= -'sd826;
        'd1456: dout <= -'sd1063;
        'd1457: dout <= -'sd1222;
        'd1458: dout <= -'sd1938;
        'd1459: dout <= -'sd1554;
        'd1460: dout <= 'sd703;
        'd1461: dout <= -'sd1241;
        'd1462: dout <= -'sd1753;
        'd1463: dout <= -'sd208;
        'd1464: dout <= -'sd876;
        'd1465: dout <= -'sd117;
        'd1466: dout <= 'sd1165;
        'd1467: dout <= -'sd1222;
        'd1468: dout <= -'sd1184;
        'd1469: dout <= 'sd1778;
        'd1470: dout <= 'sd1663;
        'd1471: dout <= -'sd956;
        'd1472: dout <= -'sd2045;
        'd1473: dout <= -'sd1652;
        'd1474: dout <= 'sd1168;
        'd1475: dout <= 'sd226;
        'd1476: dout <= 'sd19;
        'd1477: dout <= -'sd2129;
        'd1478: dout <= -'sd1606;
        'd1479: dout <= 'sd1932;
        'd1480: dout <= 'sd936;
        'd1481: dout <= -'sd148;
        'd1482: dout <= 'sd2218;
        'd1483: dout <= 'sd833;
        'd1484: dout <= 'sd1966;
        'd1485: dout <= -'sd1353;
        'd1486: dout <= -'sd1560;
        'd1487: dout <= -'sd385;
        'd1488: dout <= -'sd1280;
        'd1489: dout <= -'sd627;
        'd1490: dout <= -'sd627;
        'd1491: dout <= 'sd2099;
        'd1492: dout <= 'sd1757;
        'd1493: dout <= -'sd254;
        'd1494: dout <= -'sd602;
        'd1495: dout <= 'sd1197;
        'd1496: dout <= 'sd1436;
        'd1497: dout <= -'sd124;
        'd1498: dout <= -'sd1828;
        'd1499: dout <= 'sd1483;
        'd1500: dout <= -'sd678;
        'd1501: dout <= -'sd1235;
        'd1502: dout <= -'sd613;
        'd1503: dout <= 'sd674;
        'd1504: dout <= 'sd719;
        'd1505: dout <= 'sd1983;
        'd1506: dout <= -'sd2021;
        'd1507: dout <= 'sd1162;
        'd1508: dout <= -'sd490;
        'd1509: dout <= 'sd695;
        'd1510: dout <= 'sd1047;
        'd1511: dout <= 'sd344;
        'd1512: dout <= 'sd338;
        'd1513: dout <= -'sd818;
        'd1514: dout <= 'sd1603;
        'd1515: dout <= 'sd1864;
        'd1516: dout <= 'sd1923;
        'd1517: dout <= 'sd521;
        'd1518: dout <= -'sd145;
        'd1519: dout <= 'sd963;
        'd1520: dout <= -'sd1847;
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module hp_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [13:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'd0: dout <= 'sd1011;
        'd1: dout <= 'sd2037;
        'd2: dout <= -'sd1575;
        'd3: dout <= 'sd1189;
        'd4: dout <= 'sd2190;
        'd5: dout <= -'sd191;
        'd6: dout <= -'sd1465;
        'd7: dout <= -'sd2027;
        'd8: dout <= 'sd1501;
        'd9: dout <= 'sd1250;
        'd10: dout <= 'sd1827;
        'd11: dout <= -'sd1308;
        'd12: dout <= 'sd346;
        'd13: dout <= -'sd1585;
        'd14: dout <= -'sd2293;
        'd15: dout <= 'sd251;
        'd16: dout <= 'sd1210;
        'd17: dout <= -'sd768;
        'd18: dout <= -'sd134;
        'd19: dout <= 'sd1692;
        'd20: dout <= 'sd1681;
        'd21: dout <= -'sd1254;
        'd22: dout <= -'sd2172;
        'd23: dout <= -'sd1912;
        'd24: dout <= -'sd387;
        'd25: dout <= -'sd1544;
        'd26: dout <= 'sd1277;
        'd27: dout <= 'sd1685;
        'd28: dout <= 'sd2280;
        'd29: dout <= 'sd2005;
        'd30: dout <= -'sd1655;
        'd31: dout <= 'sd1444;
        'd32: dout <= -'sd531;
        'd33: dout <= 'sd1972;
        'd34: dout <= 'sd2210;
        'd35: dout <= 'sd445;
        'd36: dout <= -'sd1946;
        'd37: dout <= -'sd2175;
        'd38: dout <= -'sd1640;
        'd39: dout <= 'sd440;
        'd40: dout <= -'sd143;
        'd41: dout <= 'sd299;
        'd42: dout <= -'sd1570;
        'd43: dout <= -'sd76;
        'd44: dout <= 'sd1627;
        'd45: dout <= 'sd2295;
        'd46: dout <= -'sd1154;
        'd47: dout <= -'sd549;
        'd48: dout <= -'sd1575;
        'd49: dout <= 'sd507;
        'd50: dout <= -'sd1139;
        'd51: dout <= 'sd988;
        'd52: dout <= 'sd2078;
        'd53: dout <= -'sd1184;
        'd54: dout <= -'sd1486;
        'd55: dout <= 'sd1283;
        'd56: dout <= -'sd2259;
        'd57: dout <= -'sd988;
        'd58: dout <= 'sd860;
        'd59: dout <= -'sd1225;
        'd60: dout <= 'sd1837;
        'd61: dout <= 'sd1572;
        'd62: dout <= -'sd47;
        'd63: dout <= 'sd13;
        'd64: dout <= -'sd1693;
        'd65: dout <= 'sd2026;
        'd66: dout <= 'sd1509;
        'd67: dout <= 'sd7;
        'd68: dout <= 'sd958;
        'd69: dout <= 'sd1754;
        'd70: dout <= -'sd1488;
        'd71: dout <= 'sd1522;
        'd72: dout <= -'sd243;
        'd73: dout <= 'sd2047;
        'd74: dout <= 'sd936;
        'd75: dout <= -'sd1973;
        'd76: dout <= 'sd146;
        'd77: dout <= -'sd257;
        'd78: dout <= -'sd2238;
        'd79: dout <= 'sd1932;
        'd80: dout <= 'sd841;
        'd81: dout <= 'sd2259;
        'd82: dout <= -'sd979;
        'd83: dout <= 'sd2103;
        'd84: dout <= -'sd760;
        'd85: dout <= -'sd348;
        'd86: dout <= -'sd1184;
        'd87: dout <= 'sd553;
        'd88: dout <= -'sd886;
        'd89: dout <= 'sd838;
        'd90: dout <= -'sd54;
        'd91: dout <= -'sd1864;
        'd92: dout <= -'sd234;
        'd93: dout <= 'sd299;
        'd94: dout <= -'sd1784;
        'd95: dout <= -'sd1617;
        'd96: dout <= 'sd334;
        'd97: dout <= 'sd888;
        'd98: dout <= -'sd1083;
        'd99: dout <= 'sd2110;
        'd100: dout <= -'sd606;
        'd101: dout <= -'sd1387;
        'd102: dout <= -'sd589;
        'd103: dout <= -'sd2059;
        'd104: dout <= -'sd2107;
        'd105: dout <= -'sd1978;
        'd106: dout <= 'sd808;
        'd107: dout <= -'sd1157;
        'd108: dout <= 'sd228;
        'd109: dout <= 'sd57;
        'd110: dout <= 'sd1565;
        'd111: dout <= -'sd385;
        'd112: dout <= -'sd1602;
        'd113: dout <= 'sd2123;
        'd114: dout <= 'sd1370;
        'd115: dout <= -'sd1504;
        'd116: dout <= -'sd123;
        'd117: dout <= 'sd981;
        'd118: dout <= -'sd2097;
        'd119: dout <= -'sd576;
        'd120: dout <= 'sd993;
        'd121: dout <= 'sd1040;
        'd122: dout <= -'sd440;
        'd123: dout <= 'sd1411;
        'd124: dout <= -'sd2270;
        'd125: dout <= -'sd2089;
        'd126: dout <= 'sd286;
        'd127: dout <= -'sd1446;
        'd128: dout <= 'sd2014;
        'd129: dout <= 'sd1189;
        'd130: dout <= 'sd1213;
        'd131: dout <= 'sd253;
        'd132: dout <= 'sd1507;
        'd133: dout <= -'sd549;
        'd134: dout <= -'sd1186;
        'd135: dout <= 'sd1112;
        'd136: dout <= -'sd983;
        'd137: dout <= 'sd1011;
        'd138: dout <= -'sd600;
        'd139: dout <= 'sd1156;
        'd140: dout <= -'sd2189;
        'd141: dout <= 'sd1700;
        'd142: dout <= 'sd1650;
        'd143: dout <= -'sd2239;
        'd144: dout <= -'sd1715;
        'd145: dout <= -'sd41;
        'd146: dout <= 'sd1782;
        'd147: dout <= -'sd1748;
        'd148: dout <= 'sd1222;
        'd149: dout <= -'sd1628;
        'd150: dout <= -'sd1060;
        'd151: dout <= -'sd1192;
        'd152: dout <= 'sd1807;
        'd153: dout <= 'sd360;
        'd154: dout <= 'sd843;
        'd155: dout <= -'sd585;
        'd156: dout <= 'sd1504;
        'd157: dout <= -'sd2236;
        'd158: dout <= 'sd769;
        'd159: dout <= 'sd2247;
        'd160: dout <= -'sd1044;
        'd161: dout <= -'sd1485;
        'd162: dout <= 'sd1473;
        'd163: dout <= 'sd2111;
        'd164: dout <= -'sd2029;
        'd165: dout <= 'sd1522;
        'd166: dout <= -'sd963;
        'd167: dout <= 'sd66;
        'd168: dout <= -'sd153;
        'd169: dout <= 'sd1119;
        'd170: dout <= 'sd82;
        'd171: dout <= 'sd509;
        'd172: dout <= 'sd304;
        'd173: dout <= -'sd1366;
        'd174: dout <= 'sd1552;
        'd175: dout <= 'sd1851;
        'd176: dout <= -'sd854;
        'd177: dout <= 'sd299;
        'd178: dout <= -'sd1488;
        'd179: dout <= 'sd300;
        'd180: dout <= -'sd1192;
        'd181: dout <= 'sd1136;
        'd182: dout <= -'sd659;
        'd183: dout <= 'sd403;
        'd184: dout <= -'sd1544;
        'd185: dout <= 'sd1150;
        'd186: dout <= 'sd2215;
        'd187: dout <= -'sd1135;
        'd188: dout <= 'sd1468;
        'd189: dout <= 'sd336;
        'd190: dout <= 'sd2243;
        'd191: dout <= -'sd1122;
        'd192: dout <= -'sd274;
        'd193: dout <= 'sd1169;
        'd194: dout <= 'sd533;
        'd195: dout <= 'sd398;
        'd196: dout <= -'sd1563;
        'd197: dout <= 'sd696;
        'd198: dout <= 'sd346;
        'd199: dout <= 'sd1815;
        'd200: dout <= 'sd1027;
        'd201: dout <= 'sd1158;
        'd202: dout <= 'sd1786;
        'd203: dout <= -'sd105;
        'd204: dout <= -'sd199;
        'd205: dout <= 'sd1269;
        'd206: dout <= -'sd1536;
        'd207: dout <= -'sd858;
        'd208: dout <= 'sd922;
        'd209: dout <= 'sd413;
        'd210: dout <= -'sd237;
        'd211: dout <= 'sd1747;
        'd212: dout <= -'sd1940;
        'd213: dout <= 'sd50;
        'd214: dout <= 'sd2147;
        'd215: dout <= 'sd1205;
        'd216: dout <= 'sd2243;
        'd217: dout <= 'sd2282;
        'd218: dout <= 'sd2209;
        'd219: dout <= 'sd885;
        'd220: dout <= -'sd1716;
        'd221: dout <= 'sd1056;
        'd222: dout <= -'sd8;
        'd223: dout <= -'sd1604;
        'd224: dout <= 'sd1585;
        'd225: dout <= -'sd188;
        'd226: dout <= 'sd1790;
        'd227: dout <= -'sd657;
        'd228: dout <= 'sd964;
        'd229: dout <= 'sd700;
        'd230: dout <= 'sd376;
        'd231: dout <= -'sd1052;
        'd232: dout <= 'sd1938;
        'd233: dout <= -'sd55;
        'd234: dout <= -'sd591;
        'd235: dout <= -'sd1297;
        'd236: dout <= 'sd597;
        'd237: dout <= 'sd459;
        'd238: dout <= 'sd1424;
        'd239: dout <= -'sd1291;
        'd240: dout <= -'sd520;
        'd241: dout <= 'sd1808;
        'd242: dout <= -'sd1053;
        'd243: dout <= -'sd1363;
        'd244: dout <= 'sd2207;
        'd245: dout <= 'sd1082;
        'd246: dout <= -'sd2130;
        'd247: dout <= -'sd689;
        'd248: dout <= 'sd1371;
        'd249: dout <= 'sd1928;
        'd250: dout <= 'sd889;
        'd251: dout <= 'sd1099;
        'd252: dout <= -'sd358;
        'd253: dout <= -'sd1571;
        'd254: dout <= 'sd1122;
        'd255: dout <= 'sd2114;
        'd256: dout <= -'sd7;
        'd257: dout <= 'sd482;
        'd258: dout <= -'sd13;
        'd259: dout <= -'sd1365;
        'd260: dout <= -'sd2176;
        'd261: dout <= 'sd1038;
        'd262: dout <= -'sd1364;
        'd263: dout <= -'sd1243;
        'd264: dout <= 'sd697;
        'd265: dout <= 'sd1756;
        'd266: dout <= 'sd2020;
        'd267: dout <= 'sd1894;
        'd268: dout <= 'sd1916;
        'd269: dout <= -'sd6;
        'd270: dout <= 'sd960;
        'd271: dout <= 'sd2147;
        'd272: dout <= -'sd1925;
        'd273: dout <= -'sd338;
        'd274: dout <= -'sd230;
        'd275: dout <= -'sd1919;
        'd276: dout <= -'sd1949;
        'd277: dout <= -'sd1441;
        'd278: dout <= 'sd1070;
        'd279: dout <= 'sd291;
        'd280: dout <= -'sd131;
        'd281: dout <= 'sd228;
        'd282: dout <= -'sd646;
        'd283: dout <= 'sd2118;
        'd284: dout <= 'sd1359;
        'd285: dout <= -'sd587;
        'd286: dout <= -'sd1531;
        'd287: dout <= 'sd1822;
        'd288: dout <= 'sd6;
        'd289: dout <= -'sd1520;
        'd290: dout <= 'sd229;
        'd291: dout <= -'sd1259;
        'd292: dout <= -'sd1089;
        'd293: dout <= -'sd2211;
        'd294: dout <= -'sd1217;
        'd295: dout <= 'sd1161;
        'd296: dout <= -'sd496;
        'd297: dout <= 'sd1186;
        'd298: dout <= -'sd918;
        'd299: dout <= 'sd1980;
        'd300: dout <= -'sd2253;
        'd301: dout <= 'sd783;
        'd302: dout <= -'sd1696;
        'd303: dout <= -'sd712;
        'd304: dout <= -'sd2268;
        'd305: dout <= -'sd1141;
        'd306: dout <= 'sd937;
        'd307: dout <= 'sd2138;
        'd308: dout <= 'sd1604;
        'd309: dout <= 'sd2001;
        'd310: dout <= 'sd1555;
        'd311: dout <= 'sd1035;
        'd312: dout <= -'sd2113;
        'd313: dout <= -'sd1417;
        'd314: dout <= -'sd1207;
        'd315: dout <= -'sd1385;
        'd316: dout <= -'sd1469;
        'd317: dout <= -'sd1572;
        'd318: dout <= -'sd1916;
        'd319: dout <= -'sd453;
        'd320: dout <= 'sd2196;
        'd321: dout <= 'sd1450;
        'd322: dout <= -'sd506;
        'd323: dout <= 'sd2208;
        'd324: dout <= -'sd729;
        'd325: dout <= 'sd1591;
        'd326: dout <= -'sd763;
        'd327: dout <= -'sd1526;
        'd328: dout <= 'sd621;
        'd329: dout <= -'sd870;
        'd330: dout <= 'sd766;
        'd331: dout <= -'sd1112;
        'd332: dout <= -'sd655;
        'd333: dout <= 'sd736;
        'd334: dout <= -'sd1223;
        'd335: dout <= -'sd1829;
        'd336: dout <= -'sd2127;
        'd337: dout <= 'sd376;
        'd338: dout <= -'sd180;
        'd339: dout <= -'sd275;
        'd340: dout <= 'sd1087;
        'd341: dout <= -'sd561;
        'd342: dout <= -'sd720;
        'd343: dout <= -'sd753;
        'd344: dout <= 'sd1232;
        'd345: dout <= 'sd1796;
        'd346: dout <= -'sd1105;
        'd347: dout <= 'sd1631;
        'd348: dout <= -'sd880;
        'd349: dout <= 'sd1234;
        'd350: dout <= 'sd614;
        'd351: dout <= 'sd1559;
        'd352: dout <= 'sd1262;
        'd353: dout <= 'sd1589;
        'd354: dout <= -'sd143;
        'd355: dout <= 'sd1545;
        'd356: dout <= -'sd300;
        'd357: dout <= -'sd673;
        'd358: dout <= 'sd1954;
        'd359: dout <= -'sd605;
        'd360: dout <= -'sd184;
        'd361: dout <= -'sd1931;
        'd362: dout <= -'sd1681;
        'd363: dout <= 'sd1816;
        'd364: dout <= -'sd940;
        'd365: dout <= -'sd1442;
        'd366: dout <= 'sd1136;
        'd367: dout <= -'sd2213;
        'd368: dout <= -'sd1907;
        'd369: dout <= -'sd930;
        'd370: dout <= -'sd1492;
        'd371: dout <= 'sd1629;
        'd372: dout <= -'sd1289;
        'd373: dout <= 'sd955;
        'd374: dout <= -'sd803;
        'd375: dout <= -'sd1372;
        'd376: dout <= -'sd496;
        'd377: dout <= -'sd1686;
        'd378: dout <= 'sd803;
        'd379: dout <= -'sd1202;
        'd380: dout <= -'sd2113;
        'd381: dout <= 'sd175;
        'd382: dout <= 'sd1092;
        'd383: dout <= -'sd1349;
        'd384: dout <= 'sd1720;
        'd385: dout <= -'sd1802;
        'd386: dout <= -'sd2137;
        'd387: dout <= -'sd1478;
        'd388: dout <= -'sd1247;
        'd389: dout <= -'sd873;
        'd390: dout <= 'sd1681;
        'd391: dout <= 'sd676;
        'd392: dout <= 'sd1809;
        'd393: dout <= -'sd1377;
        'd394: dout <= -'sd992;
        'd395: dout <= -'sd98;
        'd396: dout <= -'sd1677;
        'd397: dout <= -'sd866;
        'd398: dout <= 'sd82;
        'd399: dout <= 'sd524;
        'd400: dout <= 'sd1166;
        'd401: dout <= -'sd614;
        'd402: dout <= -'sd2156;
        'd403: dout <= -'sd1675;
        'd404: dout <= 'sd312;
        'd405: dout <= 'sd1754;
        'd406: dout <= 'sd1781;
        'd407: dout <= 'sd2019;
        'd408: dout <= 'sd2049;
        'd409: dout <= -'sd2192;
        'd410: dout <= -'sd557;
        'd411: dout <= 'sd559;
        'd412: dout <= 'sd245;
        'd413: dout <= -'sd1141;
        'd414: dout <= -'sd321;
        'd415: dout <= 'sd802;
        'd416: dout <= -'sd2117;
        'd417: dout <= -'sd1969;
        'd418: dout <= 'sd1076;
        'd419: dout <= 'sd1537;
        'd420: dout <= 'sd490;
        'd421: dout <= 'sd859;
        'd422: dout <= 'sd1036;
        'd423: dout <= -'sd2198;
        'd424: dout <= 'sd516;
        'd425: dout <= 'sd919;
        'd426: dout <= -'sd851;
        'd427: dout <= 'sd1347;
        'd428: dout <= 'sd1522;
        'd429: dout <= 'sd2046;
        'd430: dout <= -'sd1350;
        'd431: dout <= -'sd329;
        'd432: dout <= 'sd506;
        'd433: dout <= 'sd1105;
        'd434: dout <= 'sd260;
        'd435: dout <= 'sd431;
        'd436: dout <= -'sd750;
        'd437: dout <= -'sd163;
        'd438: dout <= -'sd1638;
        'd439: dout <= -'sd1336;
        'd440: dout <= 'sd1319;
        'd441: dout <= -'sd1591;
        'd442: dout <= 'sd2238;
        'd443: dout <= -'sd332;
        'd444: dout <= -'sd1977;
        'd445: dout <= -'sd1887;
        'd446: dout <= 'sd1804;
        'd447: dout <= -'sd1946;
        'd448: dout <= 'sd2119;
        'd449: dout <= -'sd2014;
        'd450: dout <= 'sd1495;
        'd451: dout <= 'sd448;
        'd452: dout <= -'sd1658;
        'd453: dout <= 'sd989;
        'd454: dout <= 'sd700;
        'd455: dout <= -'sd321;
        'd456: dout <= -'sd9;
        'd457: dout <= -'sd120;
        'd458: dout <= 'sd497;
        'd459: dout <= -'sd306;
        'd460: dout <= -'sd1096;
        'd461: dout <= 'sd271;
        'd462: dout <= -'sd355;
        'd463: dout <= -'sd1672;
        'd464: dout <= 'sd1337;
        'd465: dout <= -'sd2051;
        'd466: dout <= -'sd824;
        'd467: dout <= 'sd1515;
        'd468: dout <= -'sd482;
        'd469: dout <= 'sd512;
        'd470: dout <= -'sd577;
        'd471: dout <= -'sd18;
        'd472: dout <= 'sd1809;
        'd473: dout <= 'sd2223;
        'd474: dout <= -'sd1820;
        'd475: dout <= 'sd1827;
        'd476: dout <= -'sd126;
        'd477: dout <= 'sd972;
        'd478: dout <= -'sd2049;
        'd479: dout <= 'sd346;
        'd480: dout <= 'sd1233;
        'd481: dout <= -'sd741;
        'd482: dout <= 'sd1814;
        'd483: dout <= 'sd620;
        'd484: dout <= -'sd1438;
        'd485: dout <= 'sd210;
        'd486: dout <= 'sd850;
        'd487: dout <= -'sd1774;
        'd488: dout <= 'sd966;
        'd489: dout <= 'sd2152;
        'd490: dout <= 'sd2195;
        'd491: dout <= -'sd1638;
        'd492: dout <= 'sd2087;
        'd493: dout <= -'sd565;
        'd494: dout <= -'sd1202;
        'd495: dout <= 'sd1459;
        'd496: dout <= -'sd1823;
        'd497: dout <= 'sd701;
        'd498: dout <= -'sd2277;
        'd499: dout <= 'sd2037;
        'd500: dout <= 'sd1147;
        'd501: dout <= -'sd689;
        'd502: dout <= 'sd606;
        'd503: dout <= -'sd2217;
        'd504: dout <= -'sd1148;
        'd505: dout <= -'sd593;
        'd506: dout <= 'sd1887;
        'd507: dout <= 'sd1981;
        'd508: dout <= -'sd643;
        'd509: dout <= 'sd2159;
        'd510: dout <= 'sd1871;
        'd511: dout <= -'sd1730;
        'd512: dout <= -'sd1091;
        'd513: dout <= 'sd1545;
        'd514: dout <= 'sd1541;
        'd515: dout <= -'sd1255;
        'd516: dout <= -'sd580;
        'd517: dout <= 'sd1436;
        'd518: dout <= 'sd543;
        'd519: dout <= -'sd251;
        'd520: dout <= -'sd340;
        'd521: dout <= 'sd554;
        'd522: dout <= 'sd1860;
        'd523: dout <= -'sd1947;
        'd524: dout <= 'sd1012;
        'd525: dout <= -'sd548;
        'd526: dout <= 'sd695;
        'd527: dout <= -'sd891;
        'd528: dout <= 'sd930;
        'd529: dout <= 'sd1249;
        'd530: dout <= 'sd1557;
        'd531: dout <= -'sd104;
        'd532: dout <= 'sd1720;
        'd533: dout <= 'sd321;
        'd534: dout <= 'sd1580;
        'd535: dout <= 'sd713;
        'd536: dout <= -'sd89;
        'd537: dout <= -'sd631;
        'd538: dout <= 'sd1323;
        'd539: dout <= 'sd1591;
        'd540: dout <= 'sd134;
        'd541: dout <= -'sd1683;
        'd542: dout <= 'sd1771;
        'd543: dout <= -'sd492;
        'd544: dout <= -'sd929;
        'd545: dout <= 'sd455;
        'd546: dout <= -'sd416;
        'd547: dout <= -'sd583;
        'd548: dout <= 'sd845;
        'd549: dout <= -'sd1343;
        'd550: dout <= -'sd1792;
        'd551: dout <= -'sd146;
        'd552: dout <= 'sd1312;
        'd553: dout <= 'sd1689;
        'd554: dout <= -'sd348;
        'd555: dout <= 'sd1436;
        'd556: dout <= -'sd755;
        'd557: dout <= 'sd1536;
        'd558: dout <= 'sd54;
        'd559: dout <= -'sd1898;
        'd560: dout <= -'sd816;
        'd561: dout <= -'sd1021;
        'd562: dout <= 'sd1663;
        'd563: dout <= 'sd421;
        'd564: dout <= 'sd860;
        'd565: dout <= 'sd2277;
        'd566: dout <= -'sd2232;
        'd567: dout <= 'sd1496;
        'd568: dout <= -'sd769;
        'd569: dout <= -'sd1411;
        'd570: dout <= -'sd999;
        'd571: dout <= 'sd1812;
        'd572: dout <= -'sd336;
        'd573: dout <= -'sd737;
        'd574: dout <= -'sd832;
        'd575: dout <= -'sd565;
        'd576: dout <= -'sd1205;
        'd577: dout <= -'sd639;
        'd578: dout <= 'sd860;
        'd579: dout <= 'sd835;
        'd580: dout <= 'sd1101;
        'd581: dout <= 'sd1340;
        'd582: dout <= -'sd102;
        'd583: dout <= 'sd1230;
        'd584: dout <= -'sd1329;
        'd585: dout <= 'sd597;
        'd586: dout <= -'sd249;
        'd587: dout <= -'sd450;
        'd588: dout <= 'sd1509;
        'd589: dout <= -'sd423;
        'd590: dout <= 'sd1731;
        'd591: dout <= -'sd1320;
        'd592: dout <= 'sd2129;
        'd593: dout <= -'sd266;
        'd594: dout <= -'sd1289;
        'd595: dout <= 'sd1142;
        'd596: dout <= -'sd754;
        'd597: dout <= -'sd1953;
        'd598: dout <= -'sd1897;
        'd599: dout <= -'sd308;
        'd600: dout <= 'sd1031;
        'd601: dout <= -'sd1106;
        'd602: dout <= -'sd388;
        'd603: dout <= -'sd2214;
        'd604: dout <= -'sd951;
        'd605: dout <= -'sd2113;
        'd606: dout <= 'sd1045;
        'd607: dout <= 'sd581;
        'd608: dout <= -'sd377;
        'd609: dout <= 'sd1814;
        'd610: dout <= 'sd1651;
        'd611: dout <= -'sd1048;
        'd612: dout <= 'sd351;
        'd613: dout <= 'sd832;
        'd614: dout <= 'sd511;
        'd615: dout <= -'sd2249;
        'd616: dout <= -'sd1466;
        'd617: dout <= -'sd1097;
        'd618: dout <= 'sd405;
        'd619: dout <= 'sd1250;
        'd620: dout <= 'sd3;
        'd621: dout <= -'sd1761;
        'd622: dout <= -'sd1474;
        'd623: dout <= -'sd1175;
        'd624: dout <= -'sd1187;
        'd625: dout <= 'sd1845;
        'd626: dout <= -'sd1525;
        'd627: dout <= -'sd111;
        'd628: dout <= -'sd1713;
        'd629: dout <= 'sd378;
        'd630: dout <= 'sd2206;
        'd631: dout <= -'sd2006;
        'd632: dout <= 'sd668;
        'd633: dout <= -'sd2107;
        'd634: dout <= 'sd196;
        'd635: dout <= 'sd521;
        'd636: dout <= 'sd1300;
        'd637: dout <= 'sd363;
        'd638: dout <= 'sd520;
        'd639: dout <= 'sd428;
        'd640: dout <= 'sd488;
        'd641: dout <= 'sd262;
        'd642: dout <= -'sd288;
        'd643: dout <= -'sd1233;
        'd644: dout <= -'sd1942;
        'd645: dout <= -'sd336;
        'd646: dout <= -'sd269;
        'd647: dout <= 'sd1281;
        'd648: dout <= 'sd796;
        'd649: dout <= -'sd884;
        'd650: dout <= 'sd1386;
        'd651: dout <= 'sd956;
        'd652: dout <= 'sd1657;
        'd653: dout <= -'sd1278;
        'd654: dout <= 'sd2124;
        'd655: dout <= -'sd404;
        'd656: dout <= -'sd456;
        'd657: dout <= -'sd2063;
        'd658: dout <= 'sd303;
        'd659: dout <= 'sd1093;
        'd660: dout <= 'sd458;
        'd661: dout <= -'sd1550;
        'd662: dout <= 'sd1834;
        'd663: dout <= 'sd2152;
        'd664: dout <= -'sd408;
        'd665: dout <= -'sd419;
        'd666: dout <= -'sd2129;
        'd667: dout <= 'sd1277;
        'd668: dout <= 'sd1063;
        'd669: dout <= 'sd810;
        'd670: dout <= -'sd648;
        'd671: dout <= -'sd1326;
        'd672: dout <= 'sd623;
        'd673: dout <= -'sd1400;
        'd674: dout <= 'sd907;
        'd675: dout <= -'sd2162;
        'd676: dout <= 'sd424;
        'd677: dout <= -'sd321;
        'd678: dout <= -'sd901;
        'd679: dout <= 'sd1618;
        'd680: dout <= 'sd946;
        'd681: dout <= 'sd2024;
        'd682: dout <= 'sd1618;
        'd683: dout <= 'sd1667;
        'd684: dout <= -'sd1042;
        'd685: dout <= 'sd27;
        'd686: dout <= 'sd860;
        'd687: dout <= 'sd885;
        'd688: dout <= 'sd1558;
        'd689: dout <= -'sd601;
        'd690: dout <= -'sd1084;
        'd691: dout <= -'sd1842;
        'd692: dout <= 'sd940;
        'd693: dout <= 'sd2047;
        'd694: dout <= 'sd365;
        'd695: dout <= -'sd807;
        'd696: dout <= 'sd2136;
        'd697: dout <= -'sd1532;
        'd698: dout <= 'sd2242;
        'd699: dout <= -'sd310;
        'd700: dout <= -'sd224;
        'd701: dout <= -'sd1731;
        'd702: dout <= -'sd348;
        'd703: dout <= -'sd406;
        'd704: dout <= -'sd674;
        'd705: dout <= 'sd611;
        'd706: dout <= -'sd1753;
        'd707: dout <= -'sd621;
        'd708: dout <= -'sd1484;
        'd709: dout <= -'sd1250;
        'd710: dout <= -'sd775;
        'd711: dout <= 'sd699;
        'd712: dout <= -'sd1401;
        'd713: dout <= -'sd1484;
        'd714: dout <= 'sd1321;
        'd715: dout <= -'sd130;
        'd716: dout <= 'sd1210;
        'd717: dout <= 'sd1541;
        'd718: dout <= 'sd1466;
        'd719: dout <= -'sd2087;
        'd720: dout <= 'sd562;
        'd721: dout <= 'sd629;
        'd722: dout <= -'sd1014;
        'd723: dout <= 'sd685;
        'd724: dout <= -'sd2156;
        'd725: dout <= -'sd194;
        'd726: dout <= -'sd1657;
        'd727: dout <= 'sd1934;
        'd728: dout <= -'sd242;
        'd729: dout <= -'sd684;
        'd730: dout <= 'sd1879;
        'd731: dout <= -'sd1279;
        'd732: dout <= 'sd1038;
        'd733: dout <= -'sd876;
        'd734: dout <= -'sd1029;
        'd735: dout <= -'sd2202;
        'd736: dout <= 'sd873;
        'd737: dout <= -'sd298;
        'd738: dout <= 'sd776;
        'd739: dout <= -'sd992;
        'd740: dout <= 'sd366;
        'd741: dout <= 'sd667;
        'd742: dout <= 'sd1823;
        'd743: dout <= -'sd324;
        'd744: dout <= -'sd890;
        'd745: dout <= -'sd712;
        'd746: dout <= -'sd1348;
        'd747: dout <= -'sd506;
        'd748: dout <= -'sd1287;
        'd749: dout <= 'sd770;
        'd750: dout <= 'sd973;
        'd751: dout <= -'sd914;
        'd752: dout <= 'sd61;
        'd753: dout <= 'sd482;
        'd754: dout <= 'sd1010;
        'd755: dout <= 'sd1923;
        'd756: dout <= 'sd38;
        'd757: dout <= 'sd1701;
        'd758: dout <= -'sd535;
        'd759: dout <= 'sd211;
        'd760: dout <= 'sd502;
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module hq1_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [13:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'd0: dout <= 'sd1237;
        'd1: dout <= 'sd153;
        'd2: dout <= -'sd2395;
        'd3: dout <= -'sd1312;
        'd4: dout <= 'sd430;
        'd5: dout <= -'sd893;
        'd6: dout <= -'sd1854;
        'd7: dout <= 'sd9;
        'd8: dout <= 'sd1221;
        'd9: dout <= 'sd3247;
        'd10: dout <= -'sd3831;
        'd11: dout <= -'sd2015;
        'd12: dout <= 'sd3706;
        'd13: dout <= -'sd3347;
        'd14: dout <= -'sd2437;
        'd15: dout <= -'sd2078;
        'd16: dout <= -'sd3738;
        'd17: dout <= 'sd968;
        'd18: dout <= -'sd3768;
        'd19: dout <= 'sd3330;
        'd20: dout <= -'sd964;
        'd21: dout <= -'sd3077;
        'd22: dout <= 'sd2115;
        'd23: dout <= 'sd2796;
        'd24: dout <= -'sd2440;
        'd25: dout <= 'sd226;
        'd26: dout <= 'sd3536;
        'd27: dout <= -'sd1097;
        'd28: dout <= 'sd3045;
        'd29: dout <= 'sd2736;
        'd30: dout <= 'sd3703;
        'd31: dout <= 'sd914;
        'd32: dout <= 'sd1174;
        'd33: dout <= 'sd409;
        'd34: dout <= -'sd2241;
        'd35: dout <= 'sd1480;
        'd36: dout <= -'sd2306;
        'd37: dout <= 'sd515;
        'd38: dout <= -'sd2855;
        'd39: dout <= -'sd3228;
        'd40: dout <= -'sd3606;
        'd41: dout <= 'sd1588;
        'd42: dout <= -'sd3644;
        'd43: dout <= -'sd1543;
        'd44: dout <= -'sd1645;
        'd45: dout <= -'sd1552;
        'd46: dout <= -'sd1198;
        'd47: dout <= -'sd214;
        'd48: dout <= 'sd1340;
        'd49: dout <= -'sd235;
        'd50: dout <= -'sd2743;
        'd51: dout <= 'sd2467;
        'd52: dout <= 'sd896;
        'd53: dout <= 'sd471;
        'd54: dout <= -'sd658;
        'd55: dout <= 'sd3119;
        'd56: dout <= -'sd355;
        'd57: dout <= -'sd2601;
        'd58: dout <= -'sd3621;
        'd59: dout <= -'sd1834;
        'd60: dout <= -'sd579;
        'd61: dout <= -'sd100;
        'd62: dout <= 'sd891;
        'd63: dout <= -'sd1300;
        'd64: dout <= 'sd3319;
        'd65: dout <= -'sd799;
        'd66: dout <= 'sd3658;
        'd67: dout <= 'sd337;
        'd68: dout <= -'sd793;
        'd69: dout <= -'sd3119;
        'd70: dout <= -'sd1250;
        'd71: dout <= -'sd2928;
        'd72: dout <= 'sd1595;
        'd73: dout <= 'sd1796;
        'd74: dout <= 'sd3714;
        'd75: dout <= 'sd2691;
        'd76: dout <= -'sd117;
        'd77: dout <= -'sd1039;
        'd78: dout <= 'sd1462;
        'd79: dout <= 'sd651;
        'd80: dout <= 'sd3182;
        'd81: dout <= 'sd274;
        'd82: dout <= -'sd2854;
        'd83: dout <= -'sd218;
        'd84: dout <= -'sd2131;
        'd85: dout <= -'sd2818;
        'd86: dout <= 'sd193;
        'd87: dout <= -'sd3352;
        'd88: dout <= -'sd894;
        'd89: dout <= -'sd3338;
        'd90: dout <= 'sd2669;
        'd91: dout <= -'sd3068;
        'd92: dout <= -'sd1244;
        'd93: dout <= 'sd501;
        'd94: dout <= 'sd831;
        'd95: dout <= 'sd988;
        'd96: dout <= 'sd3274;
        'd97: dout <= 'sd293;
        'd98: dout <= -'sd3468;
        'd99: dout <= -'sd1318;
        'd100: dout <= -'sd3589;
        'd101: dout <= -'sd40;
        'd102: dout <= 'sd2078;
        'd103: dout <= -'sd1135;
        'd104: dout <= -'sd424;
        'd105: dout <= -'sd492;
        'd106: dout <= 'sd477;
        'd107: dout <= 'sd1082;
        'd108: dout <= -'sd771;
        'd109: dout <= 'sd948;
        'd110: dout <= 'sd1915;
        'd111: dout <= -'sd2396;
        'd112: dout <= -'sd323;
        'd113: dout <= 'sd1760;
        'd114: dout <= -'sd3446;
        'd115: dout <= 'sd821;
        'd116: dout <= -'sd310;
        'd117: dout <= -'sd2120;
        'd118: dout <= -'sd488;
        'd119: dout <= -'sd122;
        'd120: dout <= 'sd3115;
        'd121: dout <= 'sd633;
        'd122: dout <= 'sd1873;
        'd123: dout <= -'sd103;
        'd124: dout <= -'sd2763;
        'd125: dout <= 'sd3310;
        'd126: dout <= 'sd386;
        'd127: dout <= -'sd3431;
        'd128: dout <= 'sd2224;
        'd129: dout <= -'sd3113;
        'd130: dout <= -'sd3623;
        'd131: dout <= 'sd3700;
        'd132: dout <= 'sd1011;
        'd133: dout <= -'sd2608;
        'd134: dout <= -'sd3054;
        'd135: dout <= 'sd1256;
        'd136: dout <= 'sd3047;
        'd137: dout <= 'sd2710;
        'd138: dout <= 'sd1456;
        'd139: dout <= -'sd2087;
        'd140: dout <= -'sd105;
        'd141: dout <= -'sd762;
        'd142: dout <= -'sd3379;
        'd143: dout <= 'sd3626;
        'd144: dout <= 'sd3429;
        'd145: dout <= 'sd1500;
        'd146: dout <= 'sd2594;
        'd147: dout <= -'sd607;
        'd148: dout <= 'sd299;
        'd149: dout <= -'sd3114;
        'd150: dout <= -'sd1825;
        'd151: dout <= 'sd3137;
        'd152: dout <= -'sd1230;
        'd153: dout <= -'sd930;
        'd154: dout <= 'sd218;
        'd155: dout <= 'sd3801;
        'd156: dout <= -'sd674;
        'd157: dout <= -'sd105;
        'd158: dout <= 'sd1842;
        'd159: dout <= 'sd349;
        'd160: dout <= 'sd1922;
        'd161: dout <= 'sd964;
        'd162: dout <= 'sd1143;
        'd163: dout <= 'sd2077;
        'd164: dout <= -'sd2907;
        'd165: dout <= -'sd2838;
        'd166: dout <= -'sd1455;
        'd167: dout <= -'sd446;
        'd168: dout <= -'sd2210;
        'd169: dout <= -'sd2006;
        'd170: dout <= 'sd2088;
        'd171: dout <= -'sd2102;
        'd172: dout <= 'sd1824;
        'd173: dout <= 'sd532;
        'd174: dout <= 'sd2357;
        'd175: dout <= -'sd3680;
        'd176: dout <= -'sd2516;
        'd177: dout <= -'sd1790;
        'd178: dout <= -'sd934;
        'd179: dout <= 'sd955;
        'd180: dout <= -'sd2061;
        'd181: dout <= 'sd3802;
        'd182: dout <= -'sd295;
        'd183: dout <= -'sd2540;
        'd184: dout <= -'sd3773;
        'd185: dout <= 'sd2433;
        'd186: dout <= 'sd2337;
        'd187: dout <= 'sd1418;
        'd188: dout <= -'sd2034;
        'd189: dout <= -'sd3794;
        'd190: dout <= -'sd478;
        'd191: dout <= -'sd2640;
        'd192: dout <= 'sd844;
        'd193: dout <= -'sd3455;
        'd194: dout <= -'sd1607;
        'd195: dout <= 'sd1936;
        'd196: dout <= 'sd2376;
        'd197: dout <= 'sd3285;
        'd198: dout <= 'sd3812;
        'd199: dout <= -'sd54;
        'd200: dout <= 'sd1833;
        'd201: dout <= -'sd2780;
        'd202: dout <= -'sd280;
        'd203: dout <= 'sd2469;
        'd204: dout <= -'sd1276;
        'd205: dout <= -'sd2630;
        'd206: dout <= -'sd281;
        'd207: dout <= 'sd925;
        'd208: dout <= 'sd1830;
        'd209: dout <= -'sd2603;
        'd210: dout <= -'sd1246;
        'd211: dout <= -'sd2270;
        'd212: dout <= -'sd3559;
        'd213: dout <= -'sd1901;
        'd214: dout <= 'sd1476;
        'd215: dout <= -'sd3128;
        'd216: dout <= 'sd841;
        'd217: dout <= -'sd3167;
        'd218: dout <= -'sd2654;
        'd219: dout <= 'sd535;
        'd220: dout <= 'sd2076;
        'd221: dout <= -'sd2516;
        'd222: dout <= 'sd3526;
        'd223: dout <= -'sd2036;
        'd224: dout <= -'sd1324;
        'd225: dout <= -'sd2787;
        'd226: dout <= -'sd3412;
        'd227: dout <= -'sd3483;
        'd228: dout <= -'sd2232;
        'd229: dout <= -'sd2644;
        'd230: dout <= 'sd3445;
        'd231: dout <= -'sd3729;
        'd232: dout <= 'sd2031;
        'd233: dout <= -'sd3830;
        'd234: dout <= -'sd3666;
        'd235: dout <= 'sd3669;
        'd236: dout <= -'sd1236;
        'd237: dout <= 'sd1723;
        'd238: dout <= -'sd1358;
        'd239: dout <= -'sd289;
        'd240: dout <= 'sd613;
        'd241: dout <= -'sd3002;
        'd242: dout <= 'sd278;
        'd243: dout <= 'sd2159;
        'd244: dout <= -'sd940;
        'd245: dout <= -'sd3055;
        'd246: dout <= -'sd3392;
        'd247: dout <= -'sd3819;
        'd248: dout <= 'sd975;
        'd249: dout <= 'sd2903;
        'd250: dout <= -'sd3145;
        'd251: dout <= 'sd2773;
        'd252: dout <= -'sd131;
        'd253: dout <= -'sd3376;
        'd254: dout <= -'sd961;
        'd255: dout <= -'sd1062;
        'd256: dout <= 'sd1212;
        'd257: dout <= 'sd833;
        'd258: dout <= -'sd1665;
        'd259: dout <= 'sd1977;
        'd260: dout <= -'sd3700;
        'd261: dout <= 'sd737;
        'd262: dout <= -'sd1697;
        'd263: dout <= -'sd1815;
        'd264: dout <= 'sd2683;
        'd265: dout <= 'sd225;
        'd266: dout <= -'sd2293;
        'd267: dout <= -'sd3188;
        'd268: dout <= 'sd3663;
        'd269: dout <= -'sd3475;
        'd270: dout <= -'sd2326;
        'd271: dout <= 'sd389;
        'd272: dout <= -'sd3192;
        'd273: dout <= 'sd2531;
        'd274: dout <= -'sd3413;
        'd275: dout <= 'sd1568;
        'd276: dout <= -'sd1500;
        'd277: dout <= -'sd1542;
        'd278: dout <= 'sd1898;
        'd279: dout <= 'sd1545;
        'd280: dout <= -'sd732;
        'd281: dout <= -'sd373;
        'd282: dout <= 'sd1411;
        'd283: dout <= -'sd529;
        'd284: dout <= -'sd1245;
        'd285: dout <= 'sd1437;
        'd286: dout <= -'sd2469;
        'd287: dout <= -'sd3794;
        'd288: dout <= -'sd2451;
        'd289: dout <= -'sd3070;
        'd290: dout <= -'sd2513;
        'd291: dout <= 'sd1004;
        'd292: dout <= 'sd2443;
        'd293: dout <= 'sd2039;
        'd294: dout <= -'sd1187;
        'd295: dout <= 'sd3444;
        'd296: dout <= 'sd77;
        'd297: dout <= -'sd1199;
        'd298: dout <= 'sd1112;
        'd299: dout <= -'sd1902;
        'd300: dout <= 'sd3628;
        'd301: dout <= -'sd255;
        'd302: dout <= 'sd918;
        'd303: dout <= 'sd3145;
        'd304: dout <= 'sd3352;
        'd305: dout <= -'sd3011;
        'd306: dout <= -'sd2152;
        'd307: dout <= 'sd3209;
        'd308: dout <= 'sd1511;
        'd309: dout <= 'sd3832;
        'd310: dout <= 'sd58;
        'd311: dout <= 'sd2658;
        'd312: dout <= 'sd1274;
        'd313: dout <= -'sd1137;
        'd314: dout <= -'sd3169;
        'd315: dout <= 'sd1219;
        'd316: dout <= -'sd2531;
        'd317: dout <= 'sd2048;
        'd318: dout <= -'sd2381;
        'd319: dout <= 'sd2163;
        'd320: dout <= -'sd1567;
        'd321: dout <= 'sd2663;
        'd322: dout <= -'sd1307;
        'd323: dout <= -'sd628;
        'd324: dout <= -'sd241;
        'd325: dout <= -'sd419;
        'd326: dout <= -'sd228;
        'd327: dout <= -'sd2494;
        'd328: dout <= -'sd72;
        'd329: dout <= 'sd2460;
        'd330: dout <= 'sd3415;
        'd331: dout <= 'sd1105;
        'd332: dout <= 'sd2348;
        'd333: dout <= -'sd3475;
        'd334: dout <= -'sd810;
        'd335: dout <= 'sd3283;
        'd336: dout <= 'sd1061;
        'd337: dout <= 'sd3803;
        'd338: dout <= -'sd899;
        'd339: dout <= 'sd2646;
        'd340: dout <= 'sd3410;
        'd341: dout <= -'sd3605;
        'd342: dout <= 'sd3335;
        'd343: dout <= -'sd1191;
        'd344: dout <= 'sd266;
        'd345: dout <= -'sd2867;
        'd346: dout <= -'sd2228;
        'd347: dout <= -'sd3596;
        'd348: dout <= -'sd409;
        'd349: dout <= -'sd2549;
        'd350: dout <= 'sd2841;
        'd351: dout <= -'sd1424;
        'd352: dout <= -'sd2418;
        'd353: dout <= -'sd3676;
        'd354: dout <= -'sd373;
        'd355: dout <= 'sd3234;
        'd356: dout <= 'sd2240;
        'd357: dout <= -'sd3235;
        'd358: dout <= 'sd2706;
        'd359: dout <= 'sd2081;
        'd360: dout <= -'sd3840;
        'd361: dout <= -'sd690;
        'd362: dout <= -'sd1882;
        'd363: dout <= -'sd1376;
        'd364: dout <= -'sd1139;
        'd365: dout <= 'sd1792;
        'd366: dout <= -'sd3711;
        'd367: dout <= -'sd140;
        'd368: dout <= -'sd3462;
        'd369: dout <= 'sd1956;
        'd370: dout <= -'sd1140;
        'd371: dout <= -'sd1346;
        'd372: dout <= 'sd898;
        'd373: dout <= -'sd1591;
        'd374: dout <= 'sd1287;
        'd375: dout <= 'sd867;
        'd376: dout <= 'sd3001;
        'd377: dout <= 'sd1039;
        'd378: dout <= -'sd800;
        'd379: dout <= -'sd1930;
        'd380: dout <= -'sd1560;
        'd381: dout <= -'sd3404;
        'd382: dout <= 'sd972;
        'd383: dout <= 'sd2140;
        'd384: dout <= 'sd3789;
        'd385: dout <= 'sd1523;
        'd386: dout <= -'sd3295;
        'd387: dout <= -'sd204;
        'd388: dout <= -'sd2745;
        'd389: dout <= -'sd159;
        'd390: dout <= -'sd3345;
        'd391: dout <= 'sd92;
        'd392: dout <= -'sd1011;
        'd393: dout <= 'sd1592;
        'd394: dout <= -'sd2388;
        'd395: dout <= 'sd1575;
        'd396: dout <= -'sd2866;
        'd397: dout <= 'sd2121;
        'd398: dout <= 'sd2325;
        'd399: dout <= 'sd2359;
        'd400: dout <= -'sd2342;
        'd401: dout <= 'sd3691;
        'd402: dout <= 'sd1152;
        'd403: dout <= 'sd2274;
        'd404: dout <= -'sd2254;
        'd405: dout <= 'sd639;
        'd406: dout <= -'sd2369;
        'd407: dout <= 'sd1064;
        'd408: dout <= 'sd533;
        'd409: dout <= -'sd3421;
        'd410: dout <= 'sd648;
        'd411: dout <= -'sd3233;
        'd412: dout <= -'sd1693;
        'd413: dout <= -'sd2899;
        'd414: dout <= 'sd2800;
        'd415: dout <= -'sd882;
        'd416: dout <= -'sd3064;
        'd417: dout <= 'sd3097;
        'd418: dout <= -'sd2122;
        'd419: dout <= -'sd2540;
        'd420: dout <= 'sd1016;
        'd421: dout <= -'sd32;
        'd422: dout <= -'sd2495;
        'd423: dout <= 'sd1140;
        'd424: dout <= 'sd707;
        'd425: dout <= -'sd3362;
        'd426: dout <= 'sd2098;
        'd427: dout <= -'sd3375;
        'd428: dout <= -'sd1586;
        'd429: dout <= -'sd2822;
        'd430: dout <= 'sd2431;
        'd431: dout <= 'sd2058;
        'd432: dout <= 'sd58;
        'd433: dout <= -'sd483;
        'd434: dout <= 'sd440;
        'd435: dout <= -'sd493;
        'd436: dout <= 'sd2891;
        'd437: dout <= -'sd3115;
        'd438: dout <= 'sd1285;
        'd439: dout <= -'sd2481;
        'd440: dout <= -'sd3790;
        'd441: dout <= 'sd2539;
        'd442: dout <= -'sd2161;
        'd443: dout <= 'sd3840;
        'd444: dout <= 'sd3398;
        'd445: dout <= -'sd1215;
        'd446: dout <= -'sd3377;
        'd447: dout <= 'sd2386;
        'd448: dout <= 'sd3661;
        'd449: dout <= 'sd1591;
        'd450: dout <= -'sd3543;
        'd451: dout <= 'sd1640;
        'd452: dout <= -'sd352;
        'd453: dout <= -'sd2544;
        'd454: dout <= -'sd858;
        'd455: dout <= -'sd2392;
        'd456: dout <= 'sd78;
        'd457: dout <= -'sd1425;
        'd458: dout <= 'sd2461;
        'd459: dout <= -'sd677;
        'd460: dout <= 'sd3671;
        'd461: dout <= 'sd671;
        'd462: dout <= 'sd1814;
        'd463: dout <= 'sd615;
        'd464: dout <= -'sd660;
        'd465: dout <= 'sd3469;
        'd466: dout <= 'sd3690;
        'd467: dout <= -'sd2523;
        'd468: dout <= 'sd3265;
        'd469: dout <= -'sd43;
        'd470: dout <= 'sd2985;
        'd471: dout <= 'sd3709;
        'd472: dout <= -'sd24;
        'd473: dout <= 'sd1246;
        'd474: dout <= -'sd1597;
        'd475: dout <= 'sd1633;
        'd476: dout <= 'sd1566;
        'd477: dout <= 'sd1781;
        'd478: dout <= 'sd3668;
        'd479: dout <= 'sd2673;
        'd480: dout <= -'sd2668;
        'd481: dout <= -'sd3651;
        'd482: dout <= -'sd2871;
        'd483: dout <= -'sd3819;
        'd484: dout <= -'sd3134;
        'd485: dout <= -'sd3302;
        'd486: dout <= 'sd3196;
        'd487: dout <= 'sd2568;
        'd488: dout <= 'sd912;
        'd489: dout <= 'sd1505;
        'd490: dout <= 'sd2074;
        'd491: dout <= 'sd629;
        'd492: dout <= 'sd3574;
        'd493: dout <= 'sd2279;
        'd494: dout <= -'sd2033;
        'd495: dout <= -'sd3705;
        'd496: dout <= -'sd605;
        'd497: dout <= 'sd1614;
        'd498: dout <= -'sd1115;
        'd499: dout <= 'sd1674;
        'd500: dout <= 'sd1020;
        'd501: dout <= 'sd2127;
        'd502: dout <= -'sd3603;
        'd503: dout <= 'sd2143;
        'd504: dout <= 'sd3508;
        'd505: dout <= -'sd3681;
        'd506: dout <= 'sd3211;
        'd507: dout <= 'sd1868;
        'd508: dout <= 'sd652;
        'd509: dout <= 'sd2982;
        'd510: dout <= 'sd2034;
        'd511: dout <= 'sd3063;
        'd512: dout <= -'sd2557;
        'd513: dout <= 'sd2477;
        'd514: dout <= -'sd1402;
        'd515: dout <= 'sd869;
        'd516: dout <= -'sd2534;
        'd517: dout <= 'sd1660;
        'd518: dout <= 'sd3348;
        'd519: dout <= -'sd1263;
        'd520: dout <= 'sd968;
        'd521: dout <= 'sd2855;
        'd522: dout <= -'sd3690;
        'd523: dout <= -'sd210;
        'd524: dout <= 'sd1231;
        'd525: dout <= -'sd171;
        'd526: dout <= -'sd888;
        'd527: dout <= -'sd202;
        'd528: dout <= 'sd1187;
        'd529: dout <= 'sd3489;
        'd530: dout <= -'sd2110;
        'd531: dout <= -'sd356;
        'd532: dout <= -'sd607;
        'd533: dout <= -'sd2774;
        'd534: dout <= 'sd3259;
        'd535: dout <= -'sd3177;
        'd536: dout <= 'sd3258;
        'd537: dout <= 'sd2789;
        'd538: dout <= -'sd3153;
        'd539: dout <= -'sd745;
        'd540: dout <= -'sd3247;
        'd541: dout <= -'sd1720;
        'd542: dout <= -'sd3189;
        'd543: dout <= 'sd3704;
        'd544: dout <= 'sd1232;
        'd545: dout <= 'sd775;
        'd546: dout <= -'sd2712;
        'd547: dout <= 'sd358;
        'd548: dout <= 'sd976;
        'd549: dout <= -'sd3154;
        'd550: dout <= -'sd1181;
        'd551: dout <= 'sd739;
        'd552: dout <= 'sd1997;
        'd553: dout <= 'sd655;
        'd554: dout <= 'sd1029;
        'd555: dout <= -'sd1882;
        'd556: dout <= 'sd701;
        'd557: dout <= -'sd2981;
        'd558: dout <= 'sd3259;
        'd559: dout <= -'sd251;
        'd560: dout <= 'sd432;
        'd561: dout <= -'sd284;
        'd562: dout <= 'sd12;
        'd563: dout <= 'sd1498;
        'd564: dout <= -'sd3399;
        'd565: dout <= 'sd213;
        'd566: dout <= -'sd2830;
        'd567: dout <= 'sd1064;
        'd568: dout <= -'sd77;
        'd569: dout <= 'sd714;
        'd570: dout <= -'sd1855;
        'd571: dout <= 'sd3588;
        'd572: dout <= 'sd3605;
        'd573: dout <= 'sd3343;
        'd574: dout <= 'sd1988;
        'd575: dout <= -'sd2424;
        'd576: dout <= -'sd3818;
        'd577: dout <= 'sd512;
        'd578: dout <= 'sd1584;
        'd579: dout <= -'sd2226;
        'd580: dout <= 'sd3458;
        'd581: dout <= -'sd679;
        'd582: dout <= 'sd652;
        'd583: dout <= -'sd3198;
        'd584: dout <= -'sd1527;
        'd585: dout <= -'sd3637;
        'd586: dout <= 'sd1654;
        'd587: dout <= 'sd2560;
        'd588: dout <= -'sd3735;
        'd589: dout <= 'sd179;
        'd590: dout <= 'sd502;
        'd591: dout <= 'sd892;
        'd592: dout <= -'sd543;
        'd593: dout <= 'sd1070;
        'd594: dout <= 'sd2251;
        'd595: dout <= -'sd2523;
        'd596: dout <= -'sd1233;
        'd597: dout <= 'sd1292;
        'd598: dout <= -'sd417;
        'd599: dout <= -'sd1244;
        'd600: dout <= 'sd1188;
        'd601: dout <= 'sd2588;
        'd602: dout <= 'sd1329;
        'd603: dout <= 'sd2078;
        'd604: dout <= -'sd172;
        'd605: dout <= -'sd2340;
        'd606: dout <= 'sd1293;
        'd607: dout <= 'sd2131;
        'd608: dout <= 'sd1652;
        'd609: dout <= -'sd3221;
        'd610: dout <= -'sd663;
        'd611: dout <= 'sd3299;
        'd612: dout <= 'sd621;
        'd613: dout <= -'sd342;
        'd614: dout <= -'sd3765;
        'd615: dout <= -'sd1718;
        'd616: dout <= -'sd454;
        'd617: dout <= -'sd1987;
        'd618: dout <= -'sd336;
        'd619: dout <= -'sd1196;
        'd620: dout <= -'sd1849;
        'd621: dout <= 'sd1578;
        'd622: dout <= -'sd2441;
        'd623: dout <= 'sd2559;
        'd624: dout <= 'sd2940;
        'd625: dout <= 'sd1133;
        'd626: dout <= 'sd1825;
        'd627: dout <= 'sd882;
        'd628: dout <= -'sd2734;
        'd629: dout <= -'sd1339;
        'd630: dout <= -'sd496;
        'd631: dout <= 'sd1211;
        'd632: dout <= -'sd399;
        'd633: dout <= -'sd1722;
        'd634: dout <= 'sd1425;
        'd635: dout <= -'sd3156;
        'd636: dout <= 'sd1312;
        'd637: dout <= 'sd3024;
        'd638: dout <= 'sd3091;
        'd639: dout <= -'sd20;
        'd640: dout <= -'sd266;
        'd641: dout <= 'sd2491;
        'd642: dout <= 'sd3546;
        'd643: dout <= -'sd3205;
        'd644: dout <= -'sd491;
        'd645: dout <= -'sd1431;
        'd646: dout <= -'sd170;
        'd647: dout <= -'sd345;
        'd648: dout <= -'sd3207;
        'd649: dout <= -'sd1269;
        'd650: dout <= -'sd1498;
        'd651: dout <= 'sd1501;
        'd652: dout <= -'sd187;
        'd653: dout <= -'sd3555;
        'd654: dout <= 'sd3608;
        'd655: dout <= -'sd2323;
        'd656: dout <= 'sd1390;
        'd657: dout <= 'sd3173;
        'd658: dout <= 'sd601;
        'd659: dout <= 'sd439;
        'd660: dout <= -'sd1508;
        'd661: dout <= 'sd2643;
        'd662: dout <= -'sd1161;
        'd663: dout <= -'sd2673;
        'd664: dout <= -'sd2319;
        'd665: dout <= -'sd2809;
        'd666: dout <= -'sd3090;
        'd667: dout <= 'sd3034;
        'd668: dout <= -'sd2342;
        'd669: dout <= 'sd2523;
        'd670: dout <= -'sd130;
        'd671: dout <= -'sd615;
        'd672: dout <= -'sd1326;
        'd673: dout <= -'sd3070;
        'd674: dout <= 'sd613;
        'd675: dout <= 'sd194;
        'd676: dout <= 'sd458;
        'd677: dout <= 'sd787;
        'd678: dout <= -'sd1107;
        'd679: dout <= -'sd26;
        'd680: dout <= 'sd2514;
        'd681: dout <= -'sd3454;
        'd682: dout <= -'sd789;
        'd683: dout <= 'sd3372;
        'd684: dout <= -'sd2227;
        'd685: dout <= -'sd1409;
        'd686: dout <= -'sd824;
        'd687: dout <= 'sd2154;
        'd688: dout <= 'sd3271;
        'd689: dout <= 'sd2025;
        'd690: dout <= 'sd1407;
        'd691: dout <= 'sd3823;
        'd692: dout <= -'sd2823;
        'd693: dout <= -'sd873;
        'd694: dout <= -'sd2328;
        'd695: dout <= 'sd3744;
        'd696: dout <= 'sd2212;
        'd697: dout <= 'sd412;
        'd698: dout <= -'sd505;
        'd699: dout <= -'sd2085;
        'd700: dout <= 'sd2473;
        'd701: dout <= 'sd3178;
        'd702: dout <= 'sd2371;
        'd703: dout <= -'sd2462;
        'd704: dout <= 'sd789;
        'd705: dout <= 'sd791;
        'd706: dout <= 'sd1956;
        'd707: dout <= -'sd3362;
        'd708: dout <= 'sd2384;
        'd709: dout <= 'sd195;
        'd710: dout <= 'sd2867;
        'd711: dout <= -'sd1699;
        'd712: dout <= -'sd1762;
        'd713: dout <= -'sd3573;
        'd714: dout <= -'sd2430;
        'd715: dout <= 'sd819;
        'd716: dout <= 'sd3439;
        'd717: dout <= 'sd1147;
        'd718: dout <= -'sd2261;
        'd719: dout <= -'sd266;
        'd720: dout <= 'sd3692;
        'd721: dout <= 'sd3699;
        'd722: dout <= -'sd1687;
        'd723: dout <= 'sd2351;
        'd724: dout <= 'sd2057;
        'd725: dout <= -'sd1917;
        'd726: dout <= 'sd3512;
        'd727: dout <= -'sd3147;
        'd728: dout <= -'sd2554;
        'd729: dout <= 'sd2700;
        'd730: dout <= 'sd2790;
        'd731: dout <= -'sd599;
        'd732: dout <= -'sd561;
        'd733: dout <= -'sd1923;
        'd734: dout <= 'sd1066;
        'd735: dout <= -'sd1798;
        'd736: dout <= -'sd3603;
        'd737: dout <= -'sd29;
        'd738: dout <= -'sd1675;
        'd739: dout <= 'sd1701;
        'd740: dout <= 'sd2822;
        'd741: dout <= 'sd3840;
        'd742: dout <= -'sd1970;
        'd743: dout <= 'sd3581;
        'd744: dout <= -'sd3792;
        'd745: dout <= 'sd1694;
        'd746: dout <= -'sd3140;
        'd747: dout <= 'sd1895;
        'd748: dout <= 'sd2734;
        'd749: dout <= 'sd2547;
        'd750: dout <= 'sd3266;
        'd751: dout <= -'sd3076;
        'd752: dout <= -'sd1468;
        'd753: dout <= -'sd1977;
        'd754: dout <= -'sd1738;
        'd755: dout <= -'sd2618;
        'd756: dout <= 'sd2039;
        'd757: dout <= 'sd3470;
        'd758: dout <= -'sd2358;
        'd759: dout <= 'sd2506;
        'd760: dout <= 'sd2121;
        'd761: dout <= -'sd1082;
        'd762: dout <= 'sd1734;
        'd763: dout <= -'sd541;
        'd764: dout <= -'sd2124;
        'd765: dout <= -'sd3695;
        'd766: dout <= -'sd1614;
        'd767: dout <= -'sd1176;
        'd768: dout <= 'sd2560;
        'd769: dout <= 'sd3415;
        'd770: dout <= -'sd1526;
        'd771: dout <= -'sd3520;
        'd772: dout <= 'sd3828;
        'd773: dout <= -'sd2040;
        'd774: dout <= 'sd2829;
        'd775: dout <= 'sd739;
        'd776: dout <= -'sd1446;
        'd777: dout <= -'sd3647;
        'd778: dout <= -'sd1082;
        'd779: dout <= 'sd1242;
        'd780: dout <= -'sd3006;
        'd781: dout <= 'sd2847;
        'd782: dout <= 'sd1548;
        'd783: dout <= 'sd625;
        'd784: dout <= 'sd1552;
        'd785: dout <= -'sd1810;
        'd786: dout <= -'sd3385;
        'd787: dout <= -'sd1995;
        'd788: dout <= -'sd1203;
        'd789: dout <= -'sd907;
        'd790: dout <= 'sd2049;
        'd791: dout <= 'sd2413;
        'd792: dout <= -'sd1723;
        'd793: dout <= -'sd2971;
        'd794: dout <= 'sd3347;
        'd795: dout <= 'sd1245;
        'd796: dout <= -'sd607;
        'd797: dout <= 'sd984;
        'd798: dout <= -'sd3135;
        'd799: dout <= 'sd280;
        'd800: dout <= 'sd1665;
        'd801: dout <= -'sd1321;
        'd802: dout <= -'sd936;
        'd803: dout <= 'sd1374;
        'd804: dout <= 'sd592;
        'd805: dout <= 'sd1134;
        'd806: dout <= 'sd2422;
        'd807: dout <= -'sd854;
        'd808: dout <= -'sd3404;
        'd809: dout <= -'sd2642;
        'd810: dout <= 'sd2389;
        'd811: dout <= -'sd3408;
        'd812: dout <= -'sd2081;
        'd813: dout <= -'sd2511;
        'd814: dout <= -'sd1897;
        'd815: dout <= 'sd1083;
        'd816: dout <= 'sd3031;
        'd817: dout <= 'sd1099;
        'd818: dout <= -'sd3173;
        'd819: dout <= -'sd519;
        'd820: dout <= -'sd788;
        'd821: dout <= 'sd1021;
        'd822: dout <= -'sd1781;
        'd823: dout <= -'sd133;
        'd824: dout <= 'sd3132;
        'd825: dout <= 'sd2397;
        'd826: dout <= 'sd1951;
        'd827: dout <= 'sd3319;
        'd828: dout <= -'sd29;
        'd829: dout <= 'sd328;
        'd830: dout <= -'sd239;
        'd831: dout <= 'sd2021;
        'd832: dout <= -'sd667;
        'd833: dout <= 'sd2093;
        'd834: dout <= -'sd3417;
        'd835: dout <= -'sd3149;
        'd836: dout <= -'sd2991;
        'd837: dout <= -'sd2550;
        'd838: dout <= -'sd669;
        'd839: dout <= 'sd1005;
        'd840: dout <= 'sd1619;
        'd841: dout <= 'sd795;
        'd842: dout <= 'sd1618;
        'd843: dout <= 'sd758;
        'd844: dout <= -'sd1098;
        'd845: dout <= 'sd3088;
        'd846: dout <= -'sd3191;
        'd847: dout <= 'sd2983;
        'd848: dout <= -'sd3531;
        'd849: dout <= 'sd3577;
        'd850: dout <= 'sd2295;
        'd851: dout <= 'sd3837;
        'd852: dout <= -'sd3468;
        'd853: dout <= 'sd184;
        'd854: dout <= -'sd1232;
        'd855: dout <= -'sd1553;
        'd856: dout <= 'sd2781;
        'd857: dout <= -'sd2447;
        'd858: dout <= -'sd1587;
        'd859: dout <= -'sd3757;
        'd860: dout <= -'sd2130;
        'd861: dout <= 'sd1616;
        'd862: dout <= -'sd1239;
        'd863: dout <= -'sd1421;
        'd864: dout <= 'sd2900;
        'd865: dout <= 'sd3674;
        'd866: dout <= 'sd2671;
        'd867: dout <= -'sd2616;
        'd868: dout <= -'sd1870;
        'd869: dout <= 'sd1173;
        'd870: dout <= -'sd3762;
        'd871: dout <= -'sd2644;
        'd872: dout <= 'sd3027;
        'd873: dout <= 'sd2752;
        'd874: dout <= 'sd2641;
        'd875: dout <= -'sd1786;
        'd876: dout <= 'sd1557;
        'd877: dout <= 'sd2756;
        'd878: dout <= 'sd2545;
        'd879: dout <= -'sd1547;
        'd880: dout <= 'sd856;
        'd881: dout <= -'sd3035;
        'd882: dout <= -'sd603;
        'd883: dout <= 'sd921;
        'd884: dout <= -'sd1581;
        'd885: dout <= 'sd1942;
        'd886: dout <= -'sd1646;
        'd887: dout <= -'sd2544;
        'd888: dout <= 'sd855;
        'd889: dout <= -'sd611;
        'd890: dout <= 'sd1074;
        'd891: dout <= -'sd943;
        'd892: dout <= -'sd2487;
        'd893: dout <= 'sd947;
        'd894: dout <= -'sd1228;
        'd895: dout <= 'sd2676;
        'd896: dout <= 'sd2221;
        'd897: dout <= -'sd1501;
        'd898: dout <= 'sd2006;
        'd899: dout <= -'sd3106;
        'd900: dout <= 'sd1003;
        'd901: dout <= 'sd162;
        'd902: dout <= 'sd2447;
        'd903: dout <= -'sd3029;
        'd904: dout <= -'sd127;
        'd905: dout <= 'sd2797;
        'd906: dout <= -'sd424;
        'd907: dout <= -'sd2480;
        'd908: dout <= -'sd3736;
        'd909: dout <= -'sd790;
        'd910: dout <= 'sd1638;
        'd911: dout <= 'sd2880;
        'd912: dout <= -'sd3106;
        'd913: dout <= 'sd1263;
        'd914: dout <= 'sd823;
        'd915: dout <= -'sd2353;
        'd916: dout <= -'sd2928;
        'd917: dout <= 'sd2953;
        'd918: dout <= -'sd2184;
        'd919: dout <= 'sd2298;
        'd920: dout <= -'sd3072;
        'd921: dout <= 'sd1656;
        'd922: dout <= 'sd1456;
        'd923: dout <= 'sd1233;
        'd924: dout <= 'sd420;
        'd925: dout <= 'sd130;
        'd926: dout <= -'sd201;
        'd927: dout <= 'sd2667;
        'd928: dout <= 'sd1840;
        'd929: dout <= -'sd2350;
        'd930: dout <= -'sd1513;
        'd931: dout <= 'sd3017;
        'd932: dout <= 'sd2266;
        'd933: dout <= -'sd426;
        'd934: dout <= 'sd783;
        'd935: dout <= -'sd1586;
        'd936: dout <= -'sd3779;
        'd937: dout <= 'sd3326;
        'd938: dout <= -'sd3158;
        'd939: dout <= -'sd1283;
        'd940: dout <= 'sd2760;
        'd941: dout <= -'sd3129;
        'd942: dout <= -'sd1690;
        'd943: dout <= -'sd3638;
        'd944: dout <= -'sd1959;
        'd945: dout <= 'sd2236;
        'd946: dout <= -'sd1011;
        'd947: dout <= 'sd3410;
        'd948: dout <= -'sd2614;
        'd949: dout <= -'sd43;
        'd950: dout <= -'sd2725;
        'd951: dout <= -'sd979;
        'd952: dout <= 'sd2666;
        'd953: dout <= 'sd2514;
        'd954: dout <= 'sd3427;
        'd955: dout <= 'sd1832;
        'd956: dout <= 'sd3599;
        'd957: dout <= 'sd2555;
        'd958: dout <= -'sd1593;
        'd959: dout <= -'sd3252;
        'd960: dout <= 'sd404;
        'd961: dout <= -'sd3730;
        'd962: dout <= -'sd2272;
        'd963: dout <= -'sd1205;
        'd964: dout <= -'sd1269;
        'd965: dout <= 'sd2402;
        'd966: dout <= -'sd1852;
        'd967: dout <= 'sd2780;
        'd968: dout <= -'sd418;
        'd969: dout <= -'sd3193;
        'd970: dout <= -'sd1126;
        'd971: dout <= -'sd1936;
        'd972: dout <= 'sd2553;
        'd973: dout <= -'sd1089;
        'd974: dout <= 'sd2486;
        'd975: dout <= -'sd1819;
        'd976: dout <= -'sd3185;
        'd977: dout <= 'sd152;
        'd978: dout <= 'sd1231;
        'd979: dout <= -'sd470;
        'd980: dout <= -'sd2308;
        'd981: dout <= -'sd691;
        'd982: dout <= -'sd61;
        'd983: dout <= -'sd1120;
        'd984: dout <= -'sd1416;
        'd985: dout <= -'sd2875;
        'd986: dout <= 'sd1816;
        'd987: dout <= 'sd1435;
        'd988: dout <= -'sd3740;
        'd989: dout <= 'sd2353;
        'd990: dout <= -'sd2154;
        'd991: dout <= 'sd629;
        'd992: dout <= -'sd1879;
        'd993: dout <= 'sd3704;
        'd994: dout <= 'sd180;
        'd995: dout <= -'sd985;
        'd996: dout <= -'sd2664;
        'd997: dout <= 'sd3217;
        'd998: dout <= 'sd2372;
        'd999: dout <= 'sd2442;
        'd1000: dout <= -'sd890;
        'd1001: dout <= -'sd190;
        'd1002: dout <= -'sd2869;
        'd1003: dout <= 'sd3548;
        'd1004: dout <= 'sd321;
        'd1005: dout <= -'sd3521;
        'd1006: dout <= -'sd474;
        'd1007: dout <= -'sd2582;
        'd1008: dout <= 'sd1665;
        'd1009: dout <= 'sd1853;
        'd1010: dout <= -'sd2368;
        'd1011: dout <= 'sd88;
        'd1012: dout <= -'sd1871;
        'd1013: dout <= -'sd2730;
        'd1014: dout <= 'sd3595;
        'd1015: dout <= -'sd3470;
        'd1016: dout <= -'sd2966;
        'd1017: dout <= -'sd3377;
        'd1018: dout <= 'sd2133;
        'd1019: dout <= -'sd1059;
        'd1020: dout <= 'sd472;
        'd1021: dout <= -'sd2521;
        'd1022: dout <= 'sd3510;
        'd1023: dout <= -'sd220;
        'd1024: dout <= 'sd632;
        'd1025: dout <= -'sd3526;
        'd1026: dout <= -'sd628;
        'd1027: dout <= -'sd1206;
        'd1028: dout <= 'sd1982;
        'd1029: dout <= 'sd3091;
        'd1030: dout <= 'sd3237;
        'd1031: dout <= 'sd3793;
        'd1032: dout <= -'sd2118;
        'd1033: dout <= 'sd3684;
        'd1034: dout <= -'sd3622;
        'd1035: dout <= -'sd617;
        'd1036: dout <= -'sd2695;
        'd1037: dout <= 'sd3105;
        'd1038: dout <= -'sd1395;
        'd1039: dout <= -'sd2834;
        'd1040: dout <= 'sd71;
        'd1041: dout <= -'sd901;
        'd1042: dout <= -'sd3443;
        'd1043: dout <= 'sd3549;
        'd1044: dout <= 'sd2863;
        'd1045: dout <= -'sd728;
        'd1046: dout <= 'sd44;
        'd1047: dout <= -'sd516;
        'd1048: dout <= -'sd123;
        'd1049: dout <= -'sd97;
        'd1050: dout <= 'sd1439;
        'd1051: dout <= -'sd1557;
        'd1052: dout <= -'sd131;
        'd1053: dout <= 'sd73;
        'd1054: dout <= -'sd191;
        'd1055: dout <= -'sd1631;
        'd1056: dout <= -'sd1262;
        'd1057: dout <= -'sd2187;
        'd1058: dout <= 'sd1505;
        'd1059: dout <= 'sd3280;
        'd1060: dout <= -'sd262;
        'd1061: dout <= 'sd855;
        'd1062: dout <= 'sd3073;
        'd1063: dout <= -'sd3639;
        'd1064: dout <= -'sd2636;
        'd1065: dout <= -'sd3045;
        'd1066: dout <= -'sd743;
        'd1067: dout <= 'sd1689;
        'd1068: dout <= 'sd2819;
        'd1069: dout <= -'sd402;
        'd1070: dout <= -'sd1762;
        'd1071: dout <= 'sd3304;
        'd1072: dout <= -'sd728;
        'd1073: dout <= 'sd3441;
        'd1074: dout <= -'sd3329;
        'd1075: dout <= 'sd1;
        'd1076: dout <= -'sd2396;
        'd1077: dout <= -'sd746;
        'd1078: dout <= 'sd2524;
        'd1079: dout <= -'sd1222;
        'd1080: dout <= -'sd2302;
        'd1081: dout <= -'sd3289;
        'd1082: dout <= -'sd3330;
        'd1083: dout <= -'sd2871;
        'd1084: dout <= 'sd119;
        'd1085: dout <= 'sd2887;
        'd1086: dout <= -'sd3531;
        'd1087: dout <= 'sd2416;
        'd1088: dout <= -'sd73;
        'd1089: dout <= -'sd520;
        'd1090: dout <= 'sd3542;
        'd1091: dout <= -'sd3728;
        'd1092: dout <= -'sd177;
        'd1093: dout <= -'sd2442;
        'd1094: dout <= -'sd125;
        'd1095: dout <= -'sd3427;
        'd1096: dout <= 'sd1731;
        'd1097: dout <= -'sd2477;
        'd1098: dout <= -'sd3328;
        'd1099: dout <= 'sd3326;
        'd1100: dout <= -'sd981;
        'd1101: dout <= 'sd2435;
        'd1102: dout <= -'sd2992;
        'd1103: dout <= 'sd557;
        'd1104: dout <= 'sd3403;
        'd1105: dout <= 'sd2203;
        'd1106: dout <= -'sd2692;
        'd1107: dout <= 'sd3811;
        'd1108: dout <= -'sd878;
        'd1109: dout <= 'sd9;
        'd1110: dout <= 'sd697;
        'd1111: dout <= 'sd3587;
        'd1112: dout <= -'sd194;
        'd1113: dout <= -'sd2010;
        'd1114: dout <= -'sd2267;
        'd1115: dout <= -'sd15;
        'd1116: dout <= -'sd2369;
        'd1117: dout <= 'sd2865;
        'd1118: dout <= 'sd2481;
        'd1119: dout <= 'sd3218;
        'd1120: dout <= 'sd3116;
        'd1121: dout <= -'sd3786;
        'd1122: dout <= -'sd1790;
        'd1123: dout <= 'sd1848;
        'd1124: dout <= 'sd1958;
        'd1125: dout <= -'sd2580;
        'd1126: dout <= -'sd2537;
        'd1127: dout <= 'sd1380;
        'd1128: dout <= -'sd83;
        'd1129: dout <= 'sd1703;
        'd1130: dout <= 'sd1748;
        'd1131: dout <= 'sd3077;
        'd1132: dout <= -'sd3203;
        'd1133: dout <= -'sd1043;
        'd1134: dout <= -'sd2585;
        'd1135: dout <= -'sd3276;
        'd1136: dout <= 'sd253;
        'd1137: dout <= -'sd1867;
        'd1138: dout <= 'sd293;
        'd1139: dout <= 'sd1114;
        'd1140: dout <= -'sd856;
        'd1141: dout <= -'sd3263;
        'd1142: dout <= -'sd745;
        'd1143: dout <= -'sd1416;
        'd1144: dout <= -'sd2683;
        'd1145: dout <= -'sd3129;
        'd1146: dout <= -'sd2919;
        'd1147: dout <= -'sd2681;
        'd1148: dout <= -'sd461;
        'd1149: dout <= -'sd3672;
        'd1150: dout <= -'sd1869;
        'd1151: dout <= -'sd3124;
        'd1152: dout <= -'sd242;
        'd1153: dout <= -'sd2326;
        'd1154: dout <= -'sd2344;
        'd1155: dout <= -'sd2299;
        'd1156: dout <= -'sd2734;
        'd1157: dout <= -'sd1359;
        'd1158: dout <= -'sd2886;
        'd1159: dout <= 'sd2000;
        'd1160: dout <= 'sd3060;
        'd1161: dout <= -'sd198;
        'd1162: dout <= 'sd99;
        'd1163: dout <= 'sd1296;
        'd1164: dout <= 'sd1652;
        'd1165: dout <= 'sd2093;
        'd1166: dout <= -'sd644;
        'd1167: dout <= -'sd2295;
        'd1168: dout <= 'sd3701;
        'd1169: dout <= -'sd2441;
        'd1170: dout <= 'sd1964;
        'd1171: dout <= -'sd618;
        'd1172: dout <= 'sd2913;
        'd1173: dout <= 'sd794;
        'd1174: dout <= -'sd3826;
        'd1175: dout <= -'sd870;
        'd1176: dout <= -'sd3378;
        'd1177: dout <= 'sd2079;
        'd1178: dout <= -'sd87;
        'd1179: dout <= -'sd2448;
        'd1180: dout <= 'sd2953;
        'd1181: dout <= 'sd2353;
        'd1182: dout <= 'sd2498;
        'd1183: dout <= -'sd262;
        'd1184: dout <= 'sd1062;
        'd1185: dout <= -'sd881;
        'd1186: dout <= -'sd2576;
        'd1187: dout <= -'sd3700;
        'd1188: dout <= 'sd2427;
        'd1189: dout <= -'sd3467;
        'd1190: dout <= 'sd2095;
        'd1191: dout <= -'sd2740;
        'd1192: dout <= 'sd452;
        'd1193: dout <= -'sd1232;
        'd1194: dout <= 'sd2980;
        'd1195: dout <= 'sd2832;
        'd1196: dout <= 'sd3627;
        'd1197: dout <= -'sd1684;
        'd1198: dout <= -'sd3693;
        'd1199: dout <= 'sd1199;
        'd1200: dout <= -'sd1157;
        'd1201: dout <= -'sd3743;
        'd1202: dout <= -'sd1051;
        'd1203: dout <= 'sd3214;
        'd1204: dout <= 'sd1094;
        'd1205: dout <= -'sd1870;
        'd1206: dout <= 'sd1369;
        'd1207: dout <= 'sd3387;
        'd1208: dout <= -'sd3553;
        'd1209: dout <= 'sd3646;
        'd1210: dout <= -'sd1528;
        'd1211: dout <= -'sd1620;
        'd1212: dout <= -'sd360;
        'd1213: dout <= 'sd1339;
        'd1214: dout <= -'sd397;
        'd1215: dout <= -'sd3806;
        'd1216: dout <= 'sd1354;
        'd1217: dout <= -'sd1220;
        'd1218: dout <= 'sd3148;
        'd1219: dout <= -'sd599;
        'd1220: dout <= -'sd3437;
        'd1221: dout <= 'sd1869;
        'd1222: dout <= 'sd3748;
        'd1223: dout <= 'sd3100;
        'd1224: dout <= 'sd1071;
        'd1225: dout <= -'sd2710;
        'd1226: dout <= -'sd2636;
        'd1227: dout <= 'sd1255;
        'd1228: dout <= -'sd137;
        'd1229: dout <= -'sd230;
        'd1230: dout <= 'sd95;
        'd1231: dout <= -'sd2920;
        'd1232: dout <= 'sd3129;
        'd1233: dout <= 'sd1895;
        'd1234: dout <= -'sd2619;
        'd1235: dout <= -'sd2694;
        'd1236: dout <= 'sd2103;
        'd1237: dout <= -'sd598;
        'd1238: dout <= 'sd1163;
        'd1239: dout <= 'sd262;
        'd1240: dout <= 'sd207;
        'd1241: dout <= -'sd2341;
        'd1242: dout <= -'sd3556;
        'd1243: dout <= 'sd1519;
        'd1244: dout <= -'sd171;
        'd1245: dout <= 'sd1640;
        'd1246: dout <= -'sd3016;
        'd1247: dout <= 'sd157;
        'd1248: dout <= -'sd2682;
        'd1249: dout <= 'sd987;
        'd1250: dout <= 'sd741;
        'd1251: dout <= -'sd370;
        'd1252: dout <= -'sd1420;
        'd1253: dout <= 'sd2673;
        'd1254: dout <= 'sd2840;
        'd1255: dout <= 'sd133;
        'd1256: dout <= -'sd2801;
        'd1257: dout <= -'sd2108;
        'd1258: dout <= -'sd626;
        'd1259: dout <= -'sd2223;
        'd1260: dout <= 'sd3647;
        'd1261: dout <= 'sd1446;
        'd1262: dout <= 'sd2085;
        'd1263: dout <= 'sd3129;
        'd1264: dout <= -'sd63;
        'd1265: dout <= -'sd603;
        'd1266: dout <= -'sd3106;
        'd1267: dout <= 'sd2281;
        'd1268: dout <= 'sd2568;
        'd1269: dout <= -'sd3714;
        'd1270: dout <= 'sd2720;
        'd1271: dout <= 'sd458;
        'd1272: dout <= 'sd3029;
        'd1273: dout <= -'sd3583;
        'd1274: dout <= -'sd1463;
        'd1275: dout <= -'sd453;
        'd1276: dout <= -'sd1917;
        'd1277: dout <= -'sd1120;
        'd1278: dout <= -'sd3170;
        'd1279: dout <= -'sd3315;
        'd1280: dout <= 'sd2580;
        'd1281: dout <= 'sd2673;
        'd1282: dout <= 'sd1983;
        'd1283: dout <= 'sd3730;
        'd1284: dout <= 'sd753;
        'd1285: dout <= -'sd3812;
        'd1286: dout <= 'sd1256;
        'd1287: dout <= 'sd1916;
        'd1288: dout <= -'sd1927;
        'd1289: dout <= -'sd1202;
        'd1290: dout <= -'sd2650;
        'd1291: dout <= 'sd3262;
        'd1292: dout <= 'sd3172;
        'd1293: dout <= -'sd77;
        'd1294: dout <= -'sd3356;
        'd1295: dout <= -'sd2795;
        'd1296: dout <= 'sd862;
        'd1297: dout <= 'sd183;
        'd1298: dout <= 'sd3836;
        'd1299: dout <= 'sd3260;
        'd1300: dout <= 'sd3820;
        'd1301: dout <= -'sd2517;
        'd1302: dout <= 'sd958;
        'd1303: dout <= -'sd2004;
        'd1304: dout <= 'sd2843;
        'd1305: dout <= 'sd2946;
        'd1306: dout <= 'sd917;
        'd1307: dout <= -'sd1837;
        'd1308: dout <= 'sd2312;
        'd1309: dout <= 'sd1228;
        'd1310: dout <= -'sd1903;
        'd1311: dout <= 'sd1092;
        'd1312: dout <= -'sd2935;
        'd1313: dout <= 'sd1737;
        'd1314: dout <= 'sd1332;
        'd1315: dout <= 'sd3119;
        'd1316: dout <= -'sd2739;
        'd1317: dout <= 'sd142;
        'd1318: dout <= 'sd1892;
        'd1319: dout <= 'sd1694;
        'd1320: dout <= 'sd2144;
        'd1321: dout <= -'sd431;
        'd1322: dout <= 'sd2220;
        'd1323: dout <= 'sd3117;
        'd1324: dout <= 'sd1282;
        'd1325: dout <= -'sd2536;
        'd1326: dout <= -'sd3733;
        'd1327: dout <= 'sd416;
        'd1328: dout <= 'sd2512;
        'd1329: dout <= -'sd1792;
        'd1330: dout <= -'sd1043;
        'd1331: dout <= -'sd1214;
        'd1332: dout <= -'sd356;
        'd1333: dout <= -'sd3772;
        'd1334: dout <= -'sd3800;
        'd1335: dout <= 'sd1907;
        'd1336: dout <= -'sd1280;
        'd1337: dout <= -'sd61;
        'd1338: dout <= 'sd1986;
        'd1339: dout <= -'sd3501;
        'd1340: dout <= 'sd2624;
        'd1341: dout <= -'sd841;
        'd1342: dout <= -'sd1;
        'd1343: dout <= -'sd668;
        'd1344: dout <= 'sd553;
        'd1345: dout <= -'sd2795;
        'd1346: dout <= 'sd1830;
        'd1347: dout <= 'sd1996;
        'd1348: dout <= 'sd2514;
        'd1349: dout <= 'sd3043;
        'd1350: dout <= -'sd3521;
        'd1351: dout <= 'sd624;
        'd1352: dout <= 'sd91;
        'd1353: dout <= 'sd2329;
        'd1354: dout <= -'sd1052;
        'd1355: dout <= 'sd624;
        'd1356: dout <= 'sd1083;
        'd1357: dout <= 'sd207;
        'd1358: dout <= -'sd1082;
        'd1359: dout <= -'sd518;
        'd1360: dout <= -'sd1070;
        'd1361: dout <= 'sd757;
        'd1362: dout <= 'sd2994;
        'd1363: dout <= 'sd3505;
        'd1364: dout <= -'sd564;
        'd1365: dout <= -'sd463;
        'd1366: dout <= 'sd2032;
        'd1367: dout <= -'sd1169;
        'd1368: dout <= -'sd2268;
        'd1369: dout <= -'sd2318;
        'd1370: dout <= 'sd2316;
        'd1371: dout <= 'sd1457;
        'd1372: dout <= 'sd3734;
        'd1373: dout <= 'sd810;
        'd1374: dout <= -'sd56;
        'd1375: dout <= -'sd2361;
        'd1376: dout <= -'sd435;
        'd1377: dout <= 'sd2698;
        'd1378: dout <= 'sd3526;
        'd1379: dout <= -'sd780;
        'd1380: dout <= 'sd1148;
        'd1381: dout <= 'sd2294;
        'd1382: dout <= -'sd614;
        'd1383: dout <= 'sd1945;
        'd1384: dout <= 'sd814;
        'd1385: dout <= -'sd2992;
        'd1386: dout <= -'sd345;
        'd1387: dout <= 'sd3736;
        'd1388: dout <= -'sd1808;
        'd1389: dout <= -'sd1620;
        'd1390: dout <= 'sd528;
        'd1391: dout <= 'sd2059;
        'd1392: dout <= -'sd3801;
        'd1393: dout <= -'sd3476;
        'd1394: dout <= -'sd720;
        'd1395: dout <= 'sd3096;
        'd1396: dout <= -'sd1170;
        'd1397: dout <= 'sd1404;
        'd1398: dout <= -'sd2571;
        'd1399: dout <= 'sd507;
        'd1400: dout <= 'sd3128;
        'd1401: dout <= 'sd2158;
        'd1402: dout <= 'sd1246;
        'd1403: dout <= 'sd2238;
        'd1404: dout <= 'sd2144;
        'd1405: dout <= -'sd286;
        'd1406: dout <= 'sd802;
        'd1407: dout <= -'sd1028;
        'd1408: dout <= 'sd394;
        'd1409: dout <= 'sd2119;
        'd1410: dout <= -'sd62;
        'd1411: dout <= 'sd514;
        'd1412: dout <= -'sd1728;
        'd1413: dout <= -'sd2411;
        'd1414: dout <= -'sd1124;
        'd1415: dout <= 'sd1351;
        'd1416: dout <= 'sd1533;
        'd1417: dout <= 'sd2721;
        'd1418: dout <= -'sd320;
        'd1419: dout <= 'sd3233;
        'd1420: dout <= 'sd866;
        'd1421: dout <= 'sd508;
        'd1422: dout <= 'sd3147;
        'd1423: dout <= 'sd1799;
        'd1424: dout <= 'sd1105;
        'd1425: dout <= 'sd3425;
        'd1426: dout <= 'sd760;
        'd1427: dout <= 'sd1048;
        'd1428: dout <= 'sd1123;
        'd1429: dout <= -'sd939;
        'd1430: dout <= -'sd307;
        'd1431: dout <= 'sd2610;
        'd1432: dout <= -'sd756;
        'd1433: dout <= -'sd2449;
        'd1434: dout <= 'sd735;
        'd1435: dout <= -'sd1621;
        'd1436: dout <= 'sd1706;
        'd1437: dout <= 'sd1887;
        'd1438: dout <= 'sd3787;
        'd1439: dout <= 'sd3644;
        'd1440: dout <= -'sd2918;
        'd1441: dout <= 'sd1375;
        'd1442: dout <= -'sd1860;
        'd1443: dout <= -'sd3792;
        'd1444: dout <= -'sd2848;
        'd1445: dout <= 'sd2708;
        'd1446: dout <= 'sd2615;
        'd1447: dout <= 'sd1592;
        'd1448: dout <= -'sd3419;
        'd1449: dout <= -'sd2880;
        'd1450: dout <= -'sd2798;
        'd1451: dout <= -'sd2682;
        'd1452: dout <= 'sd1977;
        'd1453: dout <= 'sd2899;
        'd1454: dout <= 'sd3227;
        'd1455: dout <= 'sd2224;
        'd1456: dout <= 'sd2057;
        'd1457: dout <= -'sd3159;
        'd1458: dout <= -'sd769;
        'd1459: dout <= -'sd3342;
        'd1460: dout <= 'sd2728;
        'd1461: dout <= 'sd2948;
        'd1462: dout <= -'sd1955;
        'd1463: dout <= -'sd3217;
        'd1464: dout <= -'sd1570;
        'd1465: dout <= -'sd581;
        'd1466: dout <= 'sd3423;
        'd1467: dout <= 'sd2817;
        'd1468: dout <= 'sd1684;
        'd1469: dout <= 'sd2810;
        'd1470: dout <= -'sd589;
        'd1471: dout <= 'sd3583;
        'd1472: dout <= -'sd1029;
        'd1473: dout <= -'sd392;
        'd1474: dout <= -'sd3250;
        'd1475: dout <= -'sd6;
        'd1476: dout <= 'sd2372;
        'd1477: dout <= 'sd2826;
        'd1478: dout <= -'sd3722;
        'd1479: dout <= 'sd1223;
        'd1480: dout <= -'sd14;
        'd1481: dout <= -'sd111;
        'd1482: dout <= -'sd2139;
        'd1483: dout <= -'sd988;
        'd1484: dout <= -'sd2973;
        'd1485: dout <= 'sd281;
        'd1486: dout <= 'sd2302;
        'd1487: dout <= 'sd2117;
        'd1488: dout <= -'sd2487;
        'd1489: dout <= -'sd1242;
        'd1490: dout <= -'sd1303;
        'd1491: dout <= -'sd3248;
        'd1492: dout <= 'sd2025;
        'd1493: dout <= 'sd3024;
        'd1494: dout <= 'sd3001;
        'd1495: dout <= -'sd1326;
        'd1496: dout <= -'sd523;
        'd1497: dout <= -'sd3425;
        'd1498: dout <= 'sd2959;
        'd1499: dout <= 'sd455;
        'd1500: dout <= 'sd3018;
        'd1501: dout <= -'sd2039;
        'd1502: dout <= 'sd1919;
        'd1503: dout <= -'sd2610;
        'd1504: dout <= -'sd858;
        'd1505: dout <= 'sd1610;
        'd1506: dout <= -'sd1636;
        'd1507: dout <= -'sd1186;
        'd1508: dout <= -'sd332;
        'd1509: dout <= -'sd2146;
        'd1510: dout <= -'sd1339;
        'd1511: dout <= 'sd2994;
        'd1512: dout <= 'sd3777;
        'd1513: dout <= 'sd1206;
        'd1514: dout <= 'sd784;
        'd1515: dout <= -'sd3836;
        'd1516: dout <= 'sd2021;
        'd1517: dout <= -'sd133;
        'd1518: dout <= -'sd2830;
        'd1519: dout <= 'sd694;
        'd1520: dout <= -'sd434;
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module hq2_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [13:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'd0: dout <= -'sd304;
        'd1: dout <= -'sd5981;
        'd2: dout <= -'sd854;
        'd3: dout <= -'sd2823;
        'd4: dout <= -'sd5587;
        'd5: dout <= 'sd2258;
        'd6: dout <= 'sd4430;
        'd7: dout <= 'sd4671;
        'd8: dout <= -'sd3396;
        'd9: dout <= 'sd1988;
        'd10: dout <= -'sd2194;
        'd11: dout <= -'sd867;
        'd12: dout <= -'sd2452;
        'd13: dout <= 'sd2958;
        'd14: dout <= -'sd5984;
        'd15: dout <= 'sd473;
        'd16: dout <= -'sd2029;
        'd17: dout <= -'sd516;
        'd18: dout <= -'sd2518;
        'd19: dout <= 'sd4865;
        'd20: dout <= -'sd1354;
        'd21: dout <= -'sd1707;
        'd22: dout <= 'sd5299;
        'd23: dout <= 'sd2850;
        'd24: dout <= -'sd3999;
        'd25: dout <= -'sd2172;
        'd26: dout <= -'sd742;
        'd27: dout <= -'sd5342;
        'd28: dout <= -'sd34;
        'd29: dout <= -'sd4618;
        'd30: dout <= 'sd5391;
        'd31: dout <= -'sd1880;
        'd32: dout <= -'sd3680;
        'd33: dout <= -'sd3869;
        'd34: dout <= 'sd5308;
        'd35: dout <= -'sd4834;
        'd36: dout <= -'sd5718;
        'd37: dout <= 'sd1918;
        'd38: dout <= 'sd4001;
        'd39: dout <= 'sd2510;
        'd40: dout <= -'sd3663;
        'd41: dout <= 'sd3980;
        'd42: dout <= 'sd3887;
        'd43: dout <= 'sd5473;
        'd44: dout <= 'sd5802;
        'd45: dout <= 'sd2849;
        'd46: dout <= -'sd5119;
        'd47: dout <= -'sd4396;
        'd48: dout <= -'sd5367;
        'd49: dout <= 'sd1753;
        'd50: dout <= 'sd2831;
        'd51: dout <= -'sd873;
        'd52: dout <= -'sd2339;
        'd53: dout <= -'sd2376;
        'd54: dout <= 'sd2067;
        'd55: dout <= -'sd1717;
        'd56: dout <= -'sd2936;
        'd57: dout <= 'sd724;
        'd58: dout <= 'sd2809;
        'd59: dout <= -'sd1957;
        'd60: dout <= 'sd146;
        'd61: dout <= 'sd5482;
        'd62: dout <= -'sd2074;
        'd63: dout <= -'sd3341;
        'd64: dout <= 'sd5594;
        'd65: dout <= 'sd5737;
        'd66: dout <= -'sd812;
        'd67: dout <= -'sd3237;
        'd68: dout <= 'sd2327;
        'd69: dout <= 'sd3600;
        'd70: dout <= -'sd339;
        'd71: dout <= 'sd1443;
        'd72: dout <= -'sd5030;
        'd73: dout <= 'sd4177;
        'd74: dout <= -'sd6033;
        'd75: dout <= -'sd4333;
        'd76: dout <= -'sd3649;
        'd77: dout <= 'sd2723;
        'd78: dout <= -'sd1281;
        'd79: dout <= 'sd4984;
        'd80: dout <= 'sd3562;
        'd81: dout <= 'sd4115;
        'd82: dout <= -'sd3333;
        'd83: dout <= 'sd2273;
        'd84: dout <= -'sd2913;
        'd85: dout <= 'sd1263;
        'd86: dout <= -'sd3675;
        'd87: dout <= 'sd1082;
        'd88: dout <= 'sd2992;
        'd89: dout <= -'sd1851;
        'd90: dout <= -'sd3453;
        'd91: dout <= -'sd2063;
        'd92: dout <= 'sd3694;
        'd93: dout <= 'sd3430;
        'd94: dout <= 'sd3281;
        'd95: dout <= -'sd5071;
        'd96: dout <= 'sd2775;
        'd97: dout <= -'sd3341;
        'd98: dout <= 'sd3622;
        'd99: dout <= -'sd2970;
        'd100: dout <= -'sd5284;
        'd101: dout <= -'sd5529;
        'd102: dout <= -'sd4533;
        'd103: dout <= 'sd880;
        'd104: dout <= -'sd3219;
        'd105: dout <= 'sd875;
        'd106: dout <= -'sd3421;
        'd107: dout <= 'sd4090;
        'd108: dout <= -'sd478;
        'd109: dout <= 'sd1080;
        'd110: dout <= -'sd3630;
        'd111: dout <= -'sd4785;
        'd112: dout <= 'sd5973;
        'd113: dout <= 'sd4986;
        'd114: dout <= -'sd3916;
        'd115: dout <= 'sd5033;
        'd116: dout <= -'sd2924;
        'd117: dout <= -'sd1640;
        'd118: dout <= -'sd5278;
        'd119: dout <= 'sd5682;
        'd120: dout <= 'sd1535;
        'd121: dout <= -'sd4176;
        'd122: dout <= 'sd2500;
        'd123: dout <= 'sd5656;
        'd124: dout <= -'sd461;
        'd125: dout <= 'sd5876;
        'd126: dout <= 'sd3956;
        'd127: dout <= 'sd5008;
        'd128: dout <= -'sd1301;
        'd129: dout <= -'sd2927;
        'd130: dout <= -'sd5887;
        'd131: dout <= -'sd386;
        'd132: dout <= -'sd3551;
        'd133: dout <= 'sd579;
        'd134: dout <= -'sd1876;
        'd135: dout <= -'sd3071;
        'd136: dout <= -'sd2835;
        'd137: dout <= -'sd3985;
        'd138: dout <= 'sd5386;
        'd139: dout <= 'sd5259;
        'd140: dout <= -'sd3490;
        'd141: dout <= -'sd4000;
        'd142: dout <= 'sd4352;
        'd143: dout <= -'sd4624;
        'd144: dout <= 'sd1085;
        'd145: dout <= -'sd5401;
        'd146: dout <= 'sd3089;
        'd147: dout <= -'sd2747;
        'd148: dout <= -'sd5412;
        'd149: dout <= 'sd3863;
        'd150: dout <= -'sd5294;
        'd151: dout <= 'sd1791;
        'd152: dout <= 'sd2805;
        'd153: dout <= -'sd4471;
        'd154: dout <= 'sd5417;
        'd155: dout <= -'sd4000;
        'd156: dout <= -'sd3786;
        'd157: dout <= 'sd5827;
        'd158: dout <= 'sd3632;
        'd159: dout <= -'sd5021;
        'd160: dout <= -'sd216;
        'd161: dout <= -'sd5620;
        'd162: dout <= -'sd5327;
        'd163: dout <= -'sd3893;
        'd164: dout <= 'sd5114;
        'd165: dout <= 'sd1749;
        'd166: dout <= 'sd2559;
        'd167: dout <= -'sd2808;
        'd168: dout <= 'sd4826;
        'd169: dout <= 'sd4494;
        'd170: dout <= -'sd2901;
        'd171: dout <= 'sd4497;
        'd172: dout <= 'sd4893;
        'd173: dout <= 'sd3837;
        'd174: dout <= -'sd4268;
        'd175: dout <= 'sd5993;
        'd176: dout <= 'sd1633;
        'd177: dout <= 'sd1791;
        'd178: dout <= -'sd3153;
        'd179: dout <= -'sd3991;
        'd180: dout <= 'sd5883;
        'd181: dout <= 'sd2254;
        'd182: dout <= -'sd4265;
        'd183: dout <= -'sd117;
        'd184: dout <= -'sd2665;
        'd185: dout <= -'sd4195;
        'd186: dout <= -'sd4076;
        'd187: dout <= -'sd326;
        'd188: dout <= -'sd4747;
        'd189: dout <= -'sd1518;
        'd190: dout <= 'sd5698;
        'd191: dout <= -'sd2065;
        'd192: dout <= 'sd1047;
        'd193: dout <= -'sd2579;
        'd194: dout <= -'sd4066;
        'd195: dout <= -'sd76;
        'd196: dout <= 'sd948;
        'd197: dout <= -'sd2150;
        'd198: dout <= -'sd3439;
        'd199: dout <= 'sd3063;
        'd200: dout <= -'sd1024;
        'd201: dout <= -'sd1946;
        'd202: dout <= -'sd2728;
        'd203: dout <= 'sd2118;
        'd204: dout <= -'sd1922;
        'd205: dout <= 'sd3084;
        'd206: dout <= -'sd2898;
        'd207: dout <= -'sd2564;
        'd208: dout <= -'sd5764;
        'd209: dout <= -'sd67;
        'd210: dout <= -'sd3200;
        'd211: dout <= 'sd336;
        'd212: dout <= 'sd4218;
        'd213: dout <= 'sd5943;
        'd214: dout <= 'sd5776;
        'd215: dout <= 'sd3671;
        'd216: dout <= 'sd4148;
        'd217: dout <= 'sd3862;
        'd218: dout <= 'sd5449;
        'd219: dout <= 'sd1111;
        'd220: dout <= 'sd5172;
        'd221: dout <= 'sd2092;
        'd222: dout <= 'sd1043;
        'd223: dout <= -'sd5510;
        'd224: dout <= 'sd1716;
        'd225: dout <= -'sd1948;
        'd226: dout <= 'sd2927;
        'd227: dout <= 'sd3488;
        'd228: dout <= 'sd2828;
        'd229: dout <= -'sd1388;
        'd230: dout <= 'sd2216;
        'd231: dout <= 'sd378;
        'd232: dout <= 'sd5238;
        'd233: dout <= 'sd2822;
        'd234: dout <= -'sd400;
        'd235: dout <= -'sd1307;
        'd236: dout <= 'sd2892;
        'd237: dout <= 'sd4360;
        'd238: dout <= -'sd2848;
        'd239: dout <= 'sd2005;
        'd240: dout <= -'sd3898;
        'd241: dout <= 'sd560;
        'd242: dout <= 'sd2718;
        'd243: dout <= -'sd5511;
        'd244: dout <= -'sd427;
        'd245: dout <= 'sd2012;
        'd246: dout <= -'sd186;
        'd247: dout <= -'sd1321;
        'd248: dout <= -'sd3378;
        'd249: dout <= 'sd1839;
        'd250: dout <= 'sd3133;
        'd251: dout <= 'sd1080;
        'd252: dout <= -'sd2805;
        'd253: dout <= 'sd4245;
        'd254: dout <= 'sd5992;
        'd255: dout <= 'sd3784;
        'd256: dout <= 'sd3974;
        'd257: dout <= 'sd3885;
        'd258: dout <= -'sd956;
        'd259: dout <= 'sd2752;
        'd260: dout <= -'sd1105;
        'd261: dout <= -'sd3224;
        'd262: dout <= -'sd2959;
        'd263: dout <= -'sd1824;
        'd264: dout <= -'sd2012;
        'd265: dout <= 'sd4359;
        'd266: dout <= -'sd1903;
        'd267: dout <= 'sd476;
        'd268: dout <= -'sd973;
        'd269: dout <= -'sd2282;
        'd270: dout <= 'sd393;
        'd271: dout <= 'sd536;
        'd272: dout <= 'sd10;
        'd273: dout <= -'sd1451;
        'd274: dout <= 'sd1247;
        'd275: dout <= 'sd3913;
        'd276: dout <= -'sd3238;
        'd277: dout <= -'sd1647;
        'd278: dout <= 'sd5028;
        'd279: dout <= 'sd4234;
        'd280: dout <= 'sd5004;
        'd281: dout <= -'sd3083;
        'd282: dout <= -'sd736;
        'd283: dout <= -'sd5021;
        'd284: dout <= 'sd728;
        'd285: dout <= 'sd5133;
        'd286: dout <= 'sd3747;
        'd287: dout <= -'sd5989;
        'd288: dout <= 'sd2987;
        'd289: dout <= -'sd754;
        'd290: dout <= 'sd1577;
        'd291: dout <= -'sd1598;
        'd292: dout <= 'sd2031;
        'd293: dout <= -'sd950;
        'd294: dout <= -'sd574;
        'd295: dout <= 'sd3774;
        'd296: dout <= 'sd4595;
        'd297: dout <= 'sd5391;
        'd298: dout <= -'sd1617;
        'd299: dout <= -'sd5314;
        'd300: dout <= 'sd4646;
        'd301: dout <= 'sd2827;
        'd302: dout <= 'sd5533;
        'd303: dout <= 'sd87;
        'd304: dout <= 'sd1331;
        'd305: dout <= 'sd3912;
        'd306: dout <= 'sd4754;
        'd307: dout <= -'sd6011;
        'd308: dout <= -'sd6005;
        'd309: dout <= -'sd1123;
        'd310: dout <= -'sd27;
        'd311: dout <= -'sd843;
        'd312: dout <= -'sd5585;
        'd313: dout <= -'sd4827;
        'd314: dout <= 'sd2840;
        'd315: dout <= -'sd1047;
        'd316: dout <= -'sd2648;
        'd317: dout <= 'sd4444;
        'd318: dout <= -'sd47;
        'd319: dout <= -'sd6071;
        'd320: dout <= -'sd1102;
        'd321: dout <= 'sd993;
        'd322: dout <= 'sd5193;
        'd323: dout <= -'sd5321;
        'd324: dout <= -'sd802;
        'd325: dout <= -'sd4494;
        'd326: dout <= 'sd3353;
        'd327: dout <= 'sd5438;
        'd328: dout <= 'sd5379;
        'd329: dout <= 'sd5349;
        'd330: dout <= 'sd4141;
        'd331: dout <= 'sd6101;
        'd332: dout <= 'sd1709;
        'd333: dout <= -'sd5899;
        'd334: dout <= -'sd2486;
        'd335: dout <= -'sd4321;
        'd336: dout <= -'sd3292;
        'd337: dout <= 'sd5808;
        'd338: dout <= 'sd1669;
        'd339: dout <= -'sd2711;
        'd340: dout <= 'sd217;
        'd341: dout <= -'sd5006;
        'd342: dout <= 'sd1419;
        'd343: dout <= 'sd4523;
        'd344: dout <= 'sd4627;
        'd345: dout <= 'sd2157;
        'd346: dout <= -'sd452;
        'd347: dout <= 'sd4770;
        'd348: dout <= -'sd2641;
        'd349: dout <= 'sd6074;
        'd350: dout <= 'sd3148;
        'd351: dout <= -'sd132;
        'd352: dout <= 'sd4367;
        'd353: dout <= 'sd5922;
        'd354: dout <= 'sd783;
        'd355: dout <= -'sd2620;
        'd356: dout <= -'sd1602;
        'd357: dout <= 'sd36;
        'd358: dout <= 'sd1621;
        'd359: dout <= 'sd1353;
        'd360: dout <= -'sd1271;
        'd361: dout <= -'sd331;
        'd362: dout <= -'sd556;
        'd363: dout <= 'sd4935;
        'd364: dout <= -'sd5126;
        'd365: dout <= -'sd341;
        'd366: dout <= -'sd5922;
        'd367: dout <= -'sd2765;
        'd368: dout <= 'sd4683;
        'd369: dout <= 'sd4227;
        'd370: dout <= 'sd2019;
        'd371: dout <= -'sd1016;
        'd372: dout <= 'sd4390;
        'd373: dout <= -'sd245;
        'd374: dout <= -'sd3635;
        'd375: dout <= 'sd5653;
        'd376: dout <= 'sd3689;
        'd377: dout <= -'sd2904;
        'd378: dout <= -'sd5330;
        'd379: dout <= -'sd2050;
        'd380: dout <= -'sd4167;
        'd381: dout <= -'sd916;
        'd382: dout <= 'sd1840;
        'd383: dout <= 'sd1758;
        'd384: dout <= -'sd5906;
        'd385: dout <= 'sd2034;
        'd386: dout <= 'sd4875;
        'd387: dout <= 'sd3164;
        'd388: dout <= 'sd5397;
        'd389: dout <= 'sd4579;
        'd390: dout <= -'sd4724;
        'd391: dout <= 'sd666;
        'd392: dout <= 'sd1128;
        'd393: dout <= 'sd1800;
        'd394: dout <= -'sd3904;
        'd395: dout <= -'sd5423;
        'd396: dout <= -'sd5633;
        'd397: dout <= -'sd4136;
        'd398: dout <= 'sd3927;
        'd399: dout <= 'sd2007;
        'd400: dout <= 'sd3282;
        'd401: dout <= 'sd1972;
        'd402: dout <= -'sd2639;
        'd403: dout <= -'sd5529;
        'd404: dout <= -'sd5454;
        'd405: dout <= 'sd623;
        'd406: dout <= 'sd5367;
        'd407: dout <= 'sd4437;
        'd408: dout <= 'sd2627;
        'd409: dout <= 'sd1407;
        'd410: dout <= 'sd1323;
        'd411: dout <= 'sd652;
        'd412: dout <= -'sd3764;
        'd413: dout <= -'sd3134;
        'd414: dout <= -'sd815;
        'd415: dout <= 'sd3143;
        'd416: dout <= 'sd4925;
        'd417: dout <= 'sd5512;
        'd418: dout <= -'sd2627;
        'd419: dout <= 'sd3356;
        'd420: dout <= -'sd2683;
        'd421: dout <= 'sd2055;
        'd422: dout <= 'sd1497;
        'd423: dout <= -'sd4096;
        'd424: dout <= 'sd5516;
        'd425: dout <= -'sd125;
        'd426: dout <= -'sd6060;
        'd427: dout <= 'sd509;
        'd428: dout <= 'sd6086;
        'd429: dout <= 'sd746;
        'd430: dout <= -'sd5593;
        'd431: dout <= -'sd177;
        'd432: dout <= -'sd4212;
        'd433: dout <= 'sd16;
        'd434: dout <= 'sd2765;
        'd435: dout <= -'sd4083;
        'd436: dout <= 'sd6084;
        'd437: dout <= -'sd5860;
        'd438: dout <= 'sd4322;
        'd439: dout <= -'sd3071;
        'd440: dout <= 'sd5836;
        'd441: dout <= 'sd5145;
        'd442: dout <= -'sd725;
        'd443: dout <= 'sd4188;
        'd444: dout <= -'sd1294;
        'd445: dout <= 'sd6081;
        'd446: dout <= -'sd16;
        'd447: dout <= -'sd4990;
        'd448: dout <= 'sd2055;
        'd449: dout <= -'sd5139;
        'd450: dout <= -'sd1560;
        'd451: dout <= -'sd5780;
        'd452: dout <= 'sd527;
        'd453: dout <= 'sd3123;
        'd454: dout <= 'sd5775;
        'd455: dout <= -'sd5339;
        'd456: dout <= 'sd4453;
        'd457: dout <= 'sd3474;
        'd458: dout <= 'sd5460;
        'd459: dout <= -'sd2359;
        'd460: dout <= 'sd152;
        'd461: dout <= -'sd2001;
        'd462: dout <= 'sd4512;
        'd463: dout <= 'sd407;
        'd464: dout <= -'sd2867;
        'd465: dout <= -'sd5230;
        'd466: dout <= 'sd3010;
        'd467: dout <= 'sd3406;
        'd468: dout <= 'sd4616;
        'd469: dout <= 'sd2621;
        'd470: dout <= 'sd3140;
        'd471: dout <= -'sd2452;
        'd472: dout <= 'sd3180;
        'd473: dout <= -'sd4209;
        'd474: dout <= 'sd867;
        'd475: dout <= -'sd5771;
        'd476: dout <= 'sd5782;
        'd477: dout <= -'sd1145;
        'd478: dout <= 'sd4008;
        'd479: dout <= -'sd1792;
        'd480: dout <= -'sd2323;
        'd481: dout <= -'sd2504;
        'd482: dout <= 'sd2844;
        'd483: dout <= 'sd2363;
        'd484: dout <= 'sd1504;
        'd485: dout <= -'sd3553;
        'd486: dout <= 'sd5650;
        'd487: dout <= -'sd2007;
        'd488: dout <= -'sd1816;
        'd489: dout <= 'sd3907;
        'd490: dout <= -'sd882;
        'd491: dout <= -'sd2341;
        'd492: dout <= -'sd2842;
        'd493: dout <= -'sd1358;
        'd494: dout <= 'sd2982;
        'd495: dout <= -'sd158;
        'd496: dout <= 'sd1775;
        'd497: dout <= 'sd1805;
        'd498: dout <= -'sd5497;
        'd499: dout <= 'sd2010;
        'd500: dout <= 'sd4899;
        'd501: dout <= 'sd4273;
        'd502: dout <= -'sd4828;
        'd503: dout <= 'sd4525;
        'd504: dout <= -'sd5365;
        'd505: dout <= -'sd1278;
        'd506: dout <= 'sd5841;
        'd507: dout <= 'sd2835;
        'd508: dout <= 'sd4214;
        'd509: dout <= -'sd4642;
        'd510: dout <= -'sd1235;
        'd511: dout <= -'sd2385;
        'd512: dout <= -'sd1078;
        'd513: dout <= 'sd5147;
        'd514: dout <= 'sd2930;
        'd515: dout <= -'sd3548;
        'd516: dout <= 'sd3125;
        'd517: dout <= 'sd668;
        'd518: dout <= -'sd630;
        'd519: dout <= 'sd1210;
        'd520: dout <= -'sd3307;
        'd521: dout <= -'sd3686;
        'd522: dout <= 'sd431;
        'd523: dout <= 'sd4753;
        'd524: dout <= -'sd5914;
        'd525: dout <= 'sd2675;
        'd526: dout <= -'sd5699;
        'd527: dout <= -'sd3991;
        'd528: dout <= -'sd2150;
        'd529: dout <= 'sd861;
        'd530: dout <= 'sd1015;
        'd531: dout <= 'sd5311;
        'd532: dout <= 'sd4085;
        'd533: dout <= 'sd3734;
        'd534: dout <= 'sd1853;
        'd535: dout <= -'sd2781;
        'd536: dout <= 'sd3356;
        'd537: dout <= 'sd2849;
        'd538: dout <= 'sd3522;
        'd539: dout <= 'sd2845;
        'd540: dout <= -'sd2422;
        'd541: dout <= 'sd2879;
        'd542: dout <= 'sd3736;
        'd543: dout <= 'sd2275;
        'd544: dout <= -'sd933;
        'd545: dout <= -'sd3854;
        'd546: dout <= -'sd1293;
        'd547: dout <= 'sd73;
        'd548: dout <= -'sd3291;
        'd549: dout <= -'sd1067;
        'd550: dout <= 'sd4178;
        'd551: dout <= 'sd5354;
        'd552: dout <= -'sd4942;
        'd553: dout <= -'sd3062;
        'd554: dout <= 'sd5907;
        'd555: dout <= -'sd5784;
        'd556: dout <= -'sd2808;
        'd557: dout <= 'sd3182;
        'd558: dout <= -'sd962;
        'd559: dout <= 'sd1565;
        'd560: dout <= -'sd3310;
        'd561: dout <= -'sd1217;
        'd562: dout <= -'sd1792;
        'd563: dout <= 'sd3041;
        'd564: dout <= 'sd3230;
        'd565: dout <= -'sd3708;
        'd566: dout <= -'sd5055;
        'd567: dout <= 'sd5954;
        'd568: dout <= 'sd5386;
        'd569: dout <= -'sd3107;
        'd570: dout <= -'sd5965;
        'd571: dout <= 'sd4418;
        'd572: dout <= -'sd2614;
        'd573: dout <= 'sd4717;
        'd574: dout <= 'sd3103;
        'd575: dout <= -'sd167;
        'd576: dout <= -'sd5611;
        'd577: dout <= 'sd1033;
        'd578: dout <= -'sd5442;
        'd579: dout <= 'sd2269;
        'd580: dout <= 'sd3772;
        'd581: dout <= 'sd3367;
        'd582: dout <= -'sd2801;
        'd583: dout <= -'sd1016;
        'd584: dout <= 'sd1219;
        'd585: dout <= 'sd3155;
        'd586: dout <= -'sd996;
        'd587: dout <= 'sd4922;
        'd588: dout <= 'sd5677;
        'd589: dout <= 'sd5646;
        'd590: dout <= 'sd194;
        'd591: dout <= 'sd1756;
        'd592: dout <= -'sd4749;
        'd593: dout <= -'sd6046;
        'd594: dout <= -'sd5216;
        'd595: dout <= -'sd4203;
        'd596: dout <= -'sd1677;
        'd597: dout <= -'sd798;
        'd598: dout <= -'sd441;
        'd599: dout <= -'sd596;
        'd600: dout <= -'sd3028;
        'd601: dout <= 'sd631;
        'd602: dout <= 'sd2578;
        'd603: dout <= -'sd4016;
        'd604: dout <= 'sd2994;
        'd605: dout <= 'sd805;
        'd606: dout <= -'sd2344;
        'd607: dout <= -'sd2288;
        'd608: dout <= -'sd700;
        'd609: dout <= 'sd5330;
        'd610: dout <= -'sd4446;
        'd611: dout <= 'sd4221;
        'd612: dout <= 'sd2478;
        'd613: dout <= 'sd4874;
        'd614: dout <= 'sd3781;
        'd615: dout <= 'sd43;
        'd616: dout <= 'sd3085;
        'd617: dout <= 'sd4901;
        'd618: dout <= -'sd3016;
        'd619: dout <= -'sd3578;
        'd620: dout <= 'sd677;
        'd621: dout <= -'sd3879;
        'd622: dout <= -'sd67;
        'd623: dout <= -'sd3842;
        'd624: dout <= -'sd61;
        'd625: dout <= 'sd151;
        'd626: dout <= 'sd3057;
        'd627: dout <= -'sd3943;
        'd628: dout <= 'sd3625;
        'd629: dout <= -'sd991;
        'd630: dout <= -'sd2991;
        'd631: dout <= 'sd1927;
        'd632: dout <= 'sd4044;
        'd633: dout <= 'sd6042;
        'd634: dout <= -'sd4346;
        'd635: dout <= -'sd128;
        'd636: dout <= 'sd795;
        'd637: dout <= -'sd6050;
        'd638: dout <= -'sd3737;
        'd639: dout <= 'sd2839;
        'd640: dout <= 'sd4864;
        'd641: dout <= 'sd3763;
        'd642: dout <= -'sd2956;
        'd643: dout <= -'sd3583;
        'd644: dout <= -'sd2108;
        'd645: dout <= -'sd3620;
        'd646: dout <= 'sd2580;
        'd647: dout <= -'sd1465;
        'd648: dout <= -'sd1039;
        'd649: dout <= -'sd2438;
        'd650: dout <= -'sd4387;
        'd651: dout <= 'sd4713;
        'd652: dout <= 'sd4269;
        'd653: dout <= -'sd4326;
        'd654: dout <= 'sd4902;
        'd655: dout <= -'sd2016;
        'd656: dout <= 'sd4686;
        'd657: dout <= 'sd37;
        'd658: dout <= 'sd5779;
        'd659: dout <= 'sd368;
        'd660: dout <= -'sd1774;
        'd661: dout <= -'sd4785;
        'd662: dout <= 'sd4236;
        'd663: dout <= -'sd4871;
        'd664: dout <= 'sd3816;
        'd665: dout <= 'sd5686;
        'd666: dout <= 'sd3635;
        'd667: dout <= -'sd2437;
        'd668: dout <= 'sd2810;
        'd669: dout <= 'sd5395;
        'd670: dout <= -'sd2437;
        'd671: dout <= 'sd3430;
        'd672: dout <= 'sd1181;
        'd673: dout <= 'sd4442;
        'd674: dout <= -'sd3055;
        'd675: dout <= -'sd1510;
        'd676: dout <= 'sd1430;
        'd677: dout <= -'sd3404;
        'd678: dout <= -'sd3702;
        'd679: dout <= 'sd4747;
        'd680: dout <= -'sd3409;
        'd681: dout <= -'sd393;
        'd682: dout <= -'sd2061;
        'd683: dout <= 'sd1094;
        'd684: dout <= 'sd2130;
        'd685: dout <= -'sd446;
        'd686: dout <= -'sd2075;
        'd687: dout <= -'sd2076;
        'd688: dout <= -'sd2270;
        'd689: dout <= -'sd2061;
        'd690: dout <= 'sd335;
        'd691: dout <= 'sd3475;
        'd692: dout <= -'sd2239;
        'd693: dout <= -'sd1422;
        'd694: dout <= -'sd139;
        'd695: dout <= 'sd5491;
        'd696: dout <= -'sd3092;
        'd697: dout <= 'sd5946;
        'd698: dout <= -'sd1423;
        'd699: dout <= 'sd4651;
        'd700: dout <= -'sd4707;
        'd701: dout <= -'sd2570;
        'd702: dout <= -'sd5770;
        'd703: dout <= 'sd5024;
        'd704: dout <= -'sd3708;
        'd705: dout <= -'sd5888;
        'd706: dout <= 'sd1234;
        'd707: dout <= -'sd1584;
        'd708: dout <= 'sd4450;
        'd709: dout <= 'sd1531;
        'd710: dout <= -'sd3215;
        'd711: dout <= -'sd5300;
        'd712: dout <= 'sd1694;
        'd713: dout <= 'sd4747;
        'd714: dout <= -'sd3544;
        'd715: dout <= 'sd2721;
        'd716: dout <= 'sd963;
        'd717: dout <= 'sd1386;
        'd718: dout <= 'sd2009;
        'd719: dout <= -'sd5393;
        'd720: dout <= -'sd5898;
        'd721: dout <= 'sd3271;
        'd722: dout <= 'sd1707;
        'd723: dout <= 'sd5806;
        'd724: dout <= -'sd3171;
        'd725: dout <= 'sd3681;
        'd726: dout <= -'sd6030;
        'd727: dout <= 'sd1294;
        'd728: dout <= -'sd1924;
        'd729: dout <= 'sd3935;
        'd730: dout <= 'sd430;
        'd731: dout <= -'sd628;
        'd732: dout <= 'sd2640;
        'd733: dout <= 'sd2309;
        'd734: dout <= -'sd2216;
        'd735: dout <= 'sd1226;
        'd736: dout <= -'sd6116;
        'd737: dout <= 'sd5061;
        'd738: dout <= 'sd4398;
        'd739: dout <= -'sd3568;
        'd740: dout <= -'sd384;
        'd741: dout <= 'sd1750;
        'd742: dout <= -'sd1560;
        'd743: dout <= 'sd4590;
        'd744: dout <= -'sd4572;
        'd745: dout <= -'sd910;
        'd746: dout <= -'sd3017;
        'd747: dout <= 'sd1855;
        'd748: dout <= -'sd4463;
        'd749: dout <= -'sd71;
        'd750: dout <= -'sd4482;
        'd751: dout <= 'sd4554;
        'd752: dout <= -'sd5621;
        'd753: dout <= -'sd5009;
        'd754: dout <= 'sd4085;
        'd755: dout <= -'sd2804;
        'd756: dout <= 'sd5416;
        'd757: dout <= 'sd4578;
        'd758: dout <= -'sd6092;
        'd759: dout <= -'sd2082;
        'd760: dout <= 'sd40;
        'd761: dout <= 'sd1067;
        'd762: dout <= -'sd3853;
        'd763: dout <= -'sd364;
        'd764: dout <= -'sd2476;
        'd765: dout <= 'sd3973;
        'd766: dout <= 'sd1390;
        'd767: dout <= 'sd5027;
        'd768: dout <= 'sd3178;
        'd769: dout <= -'sd3695;
        'd770: dout <= -'sd2051;
        'd771: dout <= -'sd2675;
        'd772: dout <= -'sd3853;
        'd773: dout <= -'sd808;
        'd774: dout <= 'sd2409;
        'd775: dout <= 'sd1903;
        'd776: dout <= 'sd718;
        'd777: dout <= -'sd1600;
        'd778: dout <= 'sd5408;
        'd779: dout <= -'sd3148;
        'd780: dout <= -'sd2655;
        'd781: dout <= -'sd4553;
        'd782: dout <= 'sd3015;
        'd783: dout <= -'sd6007;
        'd784: dout <= -'sd5039;
        'd785: dout <= -'sd4500;
        'd786: dout <= 'sd2304;
        'd787: dout <= 'sd2327;
        'd788: dout <= -'sd3757;
        'd789: dout <= 'sd5625;
        'd790: dout <= -'sd1478;
        'd791: dout <= 'sd1602;
        'd792: dout <= 'sd2506;
        'd793: dout <= -'sd3991;
        'd794: dout <= 'sd5764;
        'd795: dout <= 'sd728;
        'd796: dout <= -'sd4864;
        'd797: dout <= 'sd1012;
        'd798: dout <= -'sd5404;
        'd799: dout <= -'sd77;
        'd800: dout <= 'sd1589;
        'd801: dout <= 'sd2990;
        'd802: dout <= 'sd54;
        'd803: dout <= 'sd3079;
        'd804: dout <= 'sd2795;
        'd805: dout <= -'sd4269;
        'd806: dout <= 'sd91;
        'd807: dout <= -'sd4444;
        'd808: dout <= 'sd1835;
        'd809: dout <= 'sd3778;
        'd810: dout <= -'sd3755;
        'd811: dout <= -'sd672;
        'd812: dout <= 'sd3358;
        'd813: dout <= -'sd3634;
        'd814: dout <= -'sd2227;
        'd815: dout <= -'sd4012;
        'd816: dout <= 'sd3033;
        'd817: dout <= 'sd3982;
        'd818: dout <= 'sd3308;
        'd819: dout <= 'sd5813;
        'd820: dout <= -'sd3822;
        'd821: dout <= -'sd5448;
        'd822: dout <= 'sd4215;
        'd823: dout <= -'sd3024;
        'd824: dout <= -'sd1967;
        'd825: dout <= -'sd4708;
        'd826: dout <= -'sd3194;
        'd827: dout <= 'sd5423;
        'd828: dout <= -'sd4544;
        'd829: dout <= -'sd2748;
        'd830: dout <= 'sd318;
        'd831: dout <= -'sd4229;
        'd832: dout <= -'sd5432;
        'd833: dout <= -'sd1491;
        'd834: dout <= -'sd1099;
        'd835: dout <= 'sd2088;
        'd836: dout <= 'sd3316;
        'd837: dout <= 'sd1227;
        'd838: dout <= 'sd6011;
        'd839: dout <= 'sd1419;
        'd840: dout <= 'sd3116;
        'd841: dout <= 'sd3504;
        'd842: dout <= 'sd4630;
        'd843: dout <= 'sd2748;
        'd844: dout <= 'sd835;
        'd845: dout <= -'sd4548;
        'd846: dout <= 'sd3096;
        'd847: dout <= -'sd3405;
        'd848: dout <= 'sd524;
        'd849: dout <= -'sd2282;
        'd850: dout <= 'sd3005;
        'd851: dout <= 'sd3392;
        'd852: dout <= 'sd5561;
        'd853: dout <= -'sd1713;
        'd854: dout <= -'sd1246;
        'd855: dout <= -'sd4652;
        'd856: dout <= 'sd1461;
        'd857: dout <= 'sd1572;
        'd858: dout <= 'sd2647;
        'd859: dout <= 'sd3510;
        'd860: dout <= 'sd2648;
        'd861: dout <= -'sd5914;
        'd862: dout <= 'sd3831;
        'd863: dout <= -'sd1230;
        'd864: dout <= 'sd4000;
        'd865: dout <= -'sd4012;
        'd866: dout <= -'sd3694;
        'd867: dout <= -'sd1030;
        'd868: dout <= -'sd6036;
        'd869: dout <= 'sd2749;
        'd870: dout <= -'sd624;
        'd871: dout <= 'sd565;
        'd872: dout <= 'sd1367;
        'd873: dout <= 'sd5618;
        'd874: dout <= 'sd1651;
        'd875: dout <= -'sd4199;
        'd876: dout <= 'sd3244;
        'd877: dout <= -'sd4646;
        'd878: dout <= 'sd4274;
        'd879: dout <= 'sd3603;
        'd880: dout <= -'sd2944;
        'd881: dout <= 'sd3500;
        'd882: dout <= -'sd4146;
        'd883: dout <= 'sd2894;
        'd884: dout <= -'sd2748;
        'd885: dout <= 'sd1855;
        'd886: dout <= 'sd3756;
        'd887: dout <= -'sd1405;
        'd888: dout <= 'sd5765;
        'd889: dout <= -'sd2609;
        'd890: dout <= -'sd1703;
        'd891: dout <= 'sd78;
        'd892: dout <= -'sd1104;
        'd893: dout <= -'sd5085;
        'd894: dout <= 'sd676;
        'd895: dout <= -'sd1302;
        'd896: dout <= -'sd8;
        'd897: dout <= 'sd5032;
        'd898: dout <= -'sd5393;
        'd899: dout <= 'sd5362;
        'd900: dout <= 'sd1049;
        'd901: dout <= -'sd5758;
        'd902: dout <= -'sd1488;
        'd903: dout <= 'sd1486;
        'd904: dout <= -'sd1798;
        'd905: dout <= -'sd5303;
        'd906: dout <= 'sd1025;
        'd907: dout <= 'sd1640;
        'd908: dout <= 'sd1110;
        'd909: dout <= -'sd4092;
        'd910: dout <= -'sd5346;
        'd911: dout <= 'sd2543;
        'd912: dout <= -'sd4518;
        'd913: dout <= 'sd6041;
        'd914: dout <= 'sd4332;
        'd915: dout <= 'sd6040;
        'd916: dout <= -'sd495;
        'd917: dout <= 'sd930;
        'd918: dout <= -'sd2226;
        'd919: dout <= 'sd3060;
        'd920: dout <= -'sd621;
        'd921: dout <= 'sd1058;
        'd922: dout <= 'sd132;
        'd923: dout <= 'sd2627;
        'd924: dout <= 'sd2040;
        'd925: dout <= -'sd5281;
        'd926: dout <= 'sd1618;
        'd927: dout <= 'sd1036;
        'd928: dout <= 'sd754;
        'd929: dout <= 'sd2056;
        'd930: dout <= -'sd1029;
        'd931: dout <= 'sd1479;
        'd932: dout <= -'sd1380;
        'd933: dout <= 'sd5441;
        'd934: dout <= -'sd6110;
        'd935: dout <= 'sd4789;
        'd936: dout <= -'sd4025;
        'd937: dout <= 'sd4762;
        'd938: dout <= -'sd5205;
        'd939: dout <= -'sd3727;
        'd940: dout <= -'sd1717;
        'd941: dout <= 'sd415;
        'd942: dout <= 'sd313;
        'd943: dout <= 'sd1827;
        'd944: dout <= 'sd3383;
        'd945: dout <= 'sd2767;
        'd946: dout <= 'sd2657;
        'd947: dout <= -'sd1176;
        'd948: dout <= 'sd806;
        'd949: dout <= 'sd4232;
        'd950: dout <= 'sd1723;
        'd951: dout <= -'sd2970;
        'd952: dout <= 'sd2914;
        'd953: dout <= -'sd5317;
        'd954: dout <= 'sd1110;
        'd955: dout <= -'sd3900;
        'd956: dout <= 'sd2448;
        'd957: dout <= -'sd1404;
        'd958: dout <= 'sd4487;
        'd959: dout <= -'sd4890;
        'd960: dout <= 'sd2009;
        'd961: dout <= 'sd1467;
        'd962: dout <= -'sd5750;
        'd963: dout <= 'sd2200;
        'd964: dout <= -'sd4675;
        'd965: dout <= -'sd3604;
        'd966: dout <= 'sd1350;
        'd967: dout <= -'sd1316;
        'd968: dout <= -'sd2915;
        'd969: dout <= -'sd3908;
        'd970: dout <= -'sd4564;
        'd971: dout <= -'sd1217;
        'd972: dout <= -'sd259;
        'd973: dout <= 'sd5816;
        'd974: dout <= 'sd991;
        'd975: dout <= 'sd4074;
        'd976: dout <= 'sd1581;
        'd977: dout <= -'sd5300;
        'd978: dout <= 'sd1516;
        'd979: dout <= 'sd2769;
        'd980: dout <= 'sd589;
        'd981: dout <= -'sd2214;
        'd982: dout <= -'sd3482;
        'd983: dout <= -'sd4023;
        'd984: dout <= -'sd5951;
        'd985: dout <= -'sd1543;
        'd986: dout <= -'sd2040;
        'd987: dout <= -'sd4154;
        'd988: dout <= -'sd1269;
        'd989: dout <= -'sd4326;
        'd990: dout <= -'sd1368;
        'd991: dout <= -'sd2362;
        'd992: dout <= -'sd3902;
        'd993: dout <= 'sd3749;
        'd994: dout <= -'sd2702;
        'd995: dout <= 'sd3602;
        'd996: dout <= -'sd5217;
        'd997: dout <= -'sd3350;
        'd998: dout <= 'sd159;
        'd999: dout <= 'sd5806;
        'd1000: dout <= -'sd6043;
        'd1001: dout <= 'sd4357;
        'd1002: dout <= 'sd737;
        'd1003: dout <= 'sd4228;
        'd1004: dout <= 'sd4458;
        'd1005: dout <= -'sd4001;
        'd1006: dout <= -'sd966;
        'd1007: dout <= -'sd2854;
        'd1008: dout <= -'sd823;
        'd1009: dout <= -'sd425;
        'd1010: dout <= -'sd3933;
        'd1011: dout <= -'sd5650;
        'd1012: dout <= 'sd1745;
        'd1013: dout <= 'sd2127;
        'd1014: dout <= 'sd111;
        'd1015: dout <= 'sd2852;
        'd1016: dout <= -'sd3522;
        'd1017: dout <= 'sd3621;
        'd1018: dout <= 'sd5842;
        'd1019: dout <= 'sd3366;
        'd1020: dout <= -'sd870;
        'd1021: dout <= -'sd4942;
        'd1022: dout <= 'sd1478;
        'd1023: dout <= -'sd6132;
        'd1024: dout <= -'sd5989;
        'd1025: dout <= -'sd2902;
        'd1026: dout <= 'sd5391;
        'd1027: dout <= -'sd2665;
        'd1028: dout <= -'sd5256;
        'd1029: dout <= -'sd4973;
        'd1030: dout <= 'sd4545;
        'd1031: dout <= -'sd2531;
        'd1032: dout <= -'sd3601;
        'd1033: dout <= 'sd933;
        'd1034: dout <= 'sd3709;
        'd1035: dout <= -'sd5744;
        'd1036: dout <= 'sd955;
        'd1037: dout <= -'sd4356;
        'd1038: dout <= -'sd2783;
        'd1039: dout <= 'sd5653;
        'd1040: dout <= -'sd1761;
        'd1041: dout <= -'sd5883;
        'd1042: dout <= 'sd5623;
        'd1043: dout <= 'sd5330;
        'd1044: dout <= -'sd31;
        'd1045: dout <= 'sd933;
        'd1046: dout <= 'sd5501;
        'd1047: dout <= -'sd4286;
        'd1048: dout <= 'sd2478;
        'd1049: dout <= -'sd4539;
        'd1050: dout <= -'sd4768;
        'd1051: dout <= 'sd3179;
        'd1052: dout <= 'sd6122;
        'd1053: dout <= -'sd2417;
        'd1054: dout <= 'sd5696;
        'd1055: dout <= -'sd897;
        'd1056: dout <= -'sd4334;
        'd1057: dout <= 'sd2499;
        'd1058: dout <= 'sd5336;
        'd1059: dout <= 'sd1025;
        'd1060: dout <= -'sd1540;
        'd1061: dout <= -'sd3566;
        'd1062: dout <= 'sd2652;
        'd1063: dout <= 'sd975;
        'd1064: dout <= -'sd1783;
        'd1065: dout <= 'sd1275;
        'd1066: dout <= 'sd4220;
        'd1067: dout <= -'sd5771;
        'd1068: dout <= 'sd337;
        'd1069: dout <= -'sd2714;
        'd1070: dout <= -'sd2759;
        'd1071: dout <= 'sd4376;
        'd1072: dout <= -'sd4595;
        'd1073: dout <= 'sd4823;
        'd1074: dout <= 'sd5646;
        'd1075: dout <= -'sd2109;
        'd1076: dout <= -'sd5733;
        'd1077: dout <= -'sd3490;
        'd1078: dout <= 'sd4271;
        'd1079: dout <= 'sd2543;
        'd1080: dout <= -'sd2195;
        'd1081: dout <= -'sd3340;
        'd1082: dout <= -'sd3860;
        'd1083: dout <= -'sd1081;
        'd1084: dout <= -'sd5819;
        'd1085: dout <= 'sd155;
        'd1086: dout <= 'sd2010;
        'd1087: dout <= -'sd3009;
        'd1088: dout <= -'sd3733;
        'd1089: dout <= -'sd2638;
        'd1090: dout <= -'sd823;
        'd1091: dout <= 'sd2709;
        'd1092: dout <= -'sd766;
        'd1093: dout <= -'sd2471;
        'd1094: dout <= 'sd2248;
        'd1095: dout <= -'sd5983;
        'd1096: dout <= 'sd1906;
        'd1097: dout <= 'sd2961;
        'd1098: dout <= 'sd4083;
        'd1099: dout <= -'sd5333;
        'd1100: dout <= 'sd2822;
        'd1101: dout <= -'sd4925;
        'd1102: dout <= 'sd3300;
        'd1103: dout <= -'sd4573;
        'd1104: dout <= -'sd4740;
        'd1105: dout <= 'sd3236;
        'd1106: dout <= -'sd1217;
        'd1107: dout <= -'sd3031;
        'd1108: dout <= -'sd1522;
        'd1109: dout <= 'sd883;
        'd1110: dout <= -'sd5650;
        'd1111: dout <= 'sd3713;
        'd1112: dout <= -'sd384;
        'd1113: dout <= 'sd3594;
        'd1114: dout <= -'sd625;
        'd1115: dout <= -'sd3604;
        'd1116: dout <= -'sd1781;
        'd1117: dout <= 'sd1353;
        'd1118: dout <= 'sd2124;
        'd1119: dout <= -'sd1117;
        'd1120: dout <= 'sd3151;
        'd1121: dout <= 'sd788;
        'd1122: dout <= -'sd3341;
        'd1123: dout <= 'sd880;
        'd1124: dout <= -'sd3745;
        'd1125: dout <= -'sd4620;
        'd1126: dout <= -'sd384;
        'd1127: dout <= -'sd4337;
        'd1128: dout <= -'sd4289;
        'd1129: dout <= -'sd2539;
        'd1130: dout <= 'sd5840;
        'd1131: dout <= -'sd5835;
        'd1132: dout <= -'sd1470;
        'd1133: dout <= 'sd931;
        'd1134: dout <= 'sd5163;
        'd1135: dout <= -'sd3275;
        'd1136: dout <= 'sd1493;
        'd1137: dout <= -'sd1775;
        'd1138: dout <= 'sd4872;
        'd1139: dout <= -'sd2083;
        'd1140: dout <= -'sd5702;
        'd1141: dout <= -'sd4658;
        'd1142: dout <= -'sd2133;
        'd1143: dout <= 'sd670;
        'd1144: dout <= 'sd5152;
        'd1145: dout <= 'sd2859;
        'd1146: dout <= 'sd4647;
        'd1147: dout <= -'sd542;
        'd1148: dout <= -'sd1785;
        'd1149: dout <= 'sd4815;
        'd1150: dout <= 'sd221;
        'd1151: dout <= -'sd5351;
        'd1152: dout <= -'sd5809;
        'd1153: dout <= 'sd6072;
        'd1154: dout <= 'sd5538;
        'd1155: dout <= -'sd2473;
        'd1156: dout <= -'sd1223;
        'd1157: dout <= -'sd4625;
        'd1158: dout <= -'sd4678;
        'd1159: dout <= 'sd5363;
        'd1160: dout <= 'sd5167;
        'd1161: dout <= -'sd543;
        'd1162: dout <= -'sd5483;
        'd1163: dout <= 'sd3584;
        'd1164: dout <= -'sd817;
        'd1165: dout <= -'sd2869;
        'd1166: dout <= -'sd3077;
        'd1167: dout <= -'sd4759;
        'd1168: dout <= 'sd790;
        'd1169: dout <= -'sd4635;
        'd1170: dout <= 'sd3324;
        'd1171: dout <= 'sd2422;
        'd1172: dout <= -'sd1772;
        'd1173: dout <= -'sd780;
        'd1174: dout <= -'sd595;
        'd1175: dout <= -'sd6072;
        'd1176: dout <= 'sd3031;
        'd1177: dout <= -'sd4472;
        'd1178: dout <= 'sd4850;
        'd1179: dout <= -'sd4183;
        'd1180: dout <= -'sd174;
        'd1181: dout <= 'sd3186;
        'd1182: dout <= 'sd878;
        'd1183: dout <= -'sd1169;
        'd1184: dout <= 'sd5174;
        'd1185: dout <= -'sd3213;
        'd1186: dout <= -'sd975;
        'd1187: dout <= 'sd4661;
        'd1188: dout <= -'sd250;
        'd1189: dout <= 'sd602;
        'd1190: dout <= 'sd3256;
        'd1191: dout <= -'sd1366;
        'd1192: dout <= 'sd5831;
        'd1193: dout <= 'sd4338;
        'd1194: dout <= -'sd2836;
        'd1195: dout <= -'sd5005;
        'd1196: dout <= -'sd3009;
        'd1197: dout <= 'sd679;
        'd1198: dout <= 'sd1393;
        'd1199: dout <= 'sd4840;
        'd1200: dout <= 'sd3144;
        'd1201: dout <= -'sd1270;
        'd1202: dout <= -'sd6;
        'd1203: dout <= -'sd3299;
        'd1204: dout <= -'sd5834;
        'd1205: dout <= 'sd5014;
        'd1206: dout <= 'sd2714;
        'd1207: dout <= 'sd3910;
        'd1208: dout <= 'sd1828;
        'd1209: dout <= -'sd639;
        'd1210: dout <= 'sd6009;
        'd1211: dout <= 'sd716;
        'd1212: dout <= 'sd1201;
        'd1213: dout <= -'sd5035;
        'd1214: dout <= -'sd5292;
        'd1215: dout <= -'sd3777;
        'd1216: dout <= 'sd5729;
        'd1217: dout <= -'sd209;
        'd1218: dout <= -'sd5285;
        'd1219: dout <= -'sd3362;
        'd1220: dout <= -'sd1029;
        'd1221: dout <= 'sd5815;
        'd1222: dout <= -'sd2612;
        'd1223: dout <= -'sd397;
        'd1224: dout <= 'sd3979;
        'd1225: dout <= -'sd5831;
        'd1226: dout <= 'sd778;
        'd1227: dout <= 'sd4303;
        'd1228: dout <= 'sd4818;
        'd1229: dout <= 'sd4791;
        'd1230: dout <= 'sd2379;
        'd1231: dout <= 'sd1726;
        'd1232: dout <= -'sd4055;
        'd1233: dout <= 'sd786;
        'd1234: dout <= 'sd1443;
        'd1235: dout <= 'sd3692;
        'd1236: dout <= 'sd616;
        'd1237: dout <= -'sd5638;
        'd1238: dout <= -'sd927;
        'd1239: dout <= 'sd1499;
        'd1240: dout <= -'sd2638;
        'd1241: dout <= -'sd2347;
        'd1242: dout <= 'sd2539;
        'd1243: dout <= 'sd4520;
        'd1244: dout <= 'sd2084;
        'd1245: dout <= -'sd4761;
        'd1246: dout <= 'sd3855;
        'd1247: dout <= 'sd114;
        'd1248: dout <= -'sd5386;
        'd1249: dout <= 'sd2909;
        'd1250: dout <= -'sd3499;
        'd1251: dout <= -'sd4488;
        'd1252: dout <= -'sd5767;
        'd1253: dout <= 'sd4390;
        'd1254: dout <= -'sd4602;
        'd1255: dout <= -'sd3680;
        'd1256: dout <= 'sd2359;
        'd1257: dout <= 'sd5780;
        'd1258: dout <= 'sd614;
        'd1259: dout <= 'sd1676;
        'd1260: dout <= 'sd5377;
        'd1261: dout <= 'sd3444;
        'd1262: dout <= 'sd472;
        'd1263: dout <= -'sd2588;
        'd1264: dout <= -'sd4847;
        'd1265: dout <= 'sd2553;
        'd1266: dout <= -'sd291;
        'd1267: dout <= -'sd3787;
        'd1268: dout <= 'sd1719;
        'd1269: dout <= 'sd3874;
        'd1270: dout <= -'sd480;
        'd1271: dout <= 'sd2052;
        'd1272: dout <= -'sd1402;
        'd1273: dout <= -'sd1808;
        'd1274: dout <= 'sd905;
        'd1275: dout <= -'sd3431;
        'd1276: dout <= -'sd4195;
        'd1277: dout <= -'sd6061;
        'd1278: dout <= 'sd4625;
        'd1279: dout <= -'sd1381;
        'd1280: dout <= 'sd5397;
        'd1281: dout <= 'sd4742;
        'd1282: dout <= 'sd5035;
        'd1283: dout <= -'sd1801;
        'd1284: dout <= 'sd4734;
        'd1285: dout <= -'sd4281;
        'd1286: dout <= 'sd5239;
        'd1287: dout <= 'sd6001;
        'd1288: dout <= -'sd4346;
        'd1289: dout <= -'sd3971;
        'd1290: dout <= -'sd1235;
        'd1291: dout <= 'sd766;
        'd1292: dout <= 'sd2074;
        'd1293: dout <= 'sd6104;
        'd1294: dout <= 'sd2727;
        'd1295: dout <= 'sd3083;
        'd1296: dout <= -'sd1953;
        'd1297: dout <= 'sd5064;
        'd1298: dout <= 'sd3751;
        'd1299: dout <= 'sd5775;
        'd1300: dout <= -'sd1053;
        'd1301: dout <= 'sd5266;
        'd1302: dout <= -'sd1042;
        'd1303: dout <= 'sd398;
        'd1304: dout <= 'sd1218;
        'd1305: dout <= -'sd2465;
        'd1306: dout <= 'sd2215;
        'd1307: dout <= 'sd252;
        'd1308: dout <= -'sd4617;
        'd1309: dout <= -'sd3082;
        'd1310: dout <= -'sd4316;
        'd1311: dout <= -'sd2263;
        'd1312: dout <= -'sd2422;
        'd1313: dout <= 'sd4785;
        'd1314: dout <= -'sd4021;
        'd1315: dout <= -'sd5990;
        'd1316: dout <= -'sd1636;
        'd1317: dout <= 'sd2230;
        'd1318: dout <= 'sd2312;
        'd1319: dout <= 'sd673;
        'd1320: dout <= -'sd4620;
        'd1321: dout <= 'sd3718;
        'd1322: dout <= -'sd2163;
        'd1323: dout <= 'sd372;
        'd1324: dout <= 'sd6121;
        'd1325: dout <= 'sd2582;
        'd1326: dout <= 'sd1771;
        'd1327: dout <= -'sd3802;
        'd1328: dout <= -'sd5403;
        'd1329: dout <= 'sd4233;
        'd1330: dout <= -'sd5645;
        'd1331: dout <= 'sd1794;
        'd1332: dout <= 'sd5694;
        'd1333: dout <= 'sd3004;
        'd1334: dout <= 'sd1685;
        'd1335: dout <= 'sd3133;
        'd1336: dout <= 'sd4284;
        'd1337: dout <= 'sd3234;
        'd1338: dout <= -'sd481;
        'd1339: dout <= 'sd1080;
        'd1340: dout <= -'sd2899;
        'd1341: dout <= 'sd782;
        'd1342: dout <= -'sd5253;
        'd1343: dout <= -'sd4106;
        'd1344: dout <= 'sd3188;
        'd1345: dout <= 'sd1669;
        'd1346: dout <= -'sd700;
        'd1347: dout <= 'sd146;
        'd1348: dout <= 'sd3413;
        'd1349: dout <= 'sd918;
        'd1350: dout <= -'sd2433;
        'd1351: dout <= 'sd1472;
        'd1352: dout <= 'sd1345;
        'd1353: dout <= 'sd5490;
        'd1354: dout <= -'sd5261;
        'd1355: dout <= -'sd2446;
        'd1356: dout <= 'sd3706;
        'd1357: dout <= -'sd2941;
        'd1358: dout <= -'sd3;
        'd1359: dout <= 'sd3918;
        'd1360: dout <= -'sd212;
        'd1361: dout <= -'sd5207;
        'd1362: dout <= -'sd70;
        'd1363: dout <= 'sd5499;
        'd1364: dout <= -'sd383;
        'd1365: dout <= 'sd361;
        'd1366: dout <= -'sd4596;
        'd1367: dout <= 'sd3709;
        'd1368: dout <= 'sd4322;
        'd1369: dout <= 'sd4581;
        'd1370: dout <= 'sd1362;
        'd1371: dout <= -'sd3345;
        'd1372: dout <= -'sd903;
        'd1373: dout <= -'sd864;
        'd1374: dout <= 'sd723;
        'd1375: dout <= -'sd4661;
        'd1376: dout <= 'sd4487;
        'd1377: dout <= -'sd248;
        'd1378: dout <= 'sd3859;
        'd1379: dout <= 'sd2500;
        'd1380: dout <= 'sd4356;
        'd1381: dout <= 'sd2390;
        'd1382: dout <= 'sd1278;
        'd1383: dout <= 'sd2674;
        'd1384: dout <= 'sd5640;
        'd1385: dout <= 'sd5432;
        'd1386: dout <= -'sd1277;
        'd1387: dout <= 'sd4749;
        'd1388: dout <= -'sd4138;
        'd1389: dout <= 'sd6002;
        'd1390: dout <= -'sd2426;
        'd1391: dout <= -'sd5415;
        'd1392: dout <= -'sd3765;
        'd1393: dout <= -'sd4237;
        'd1394: dout <= -'sd5052;
        'd1395: dout <= 'sd1011;
        'd1396: dout <= -'sd4810;
        'd1397: dout <= -'sd3756;
        'd1398: dout <= -'sd3513;
        'd1399: dout <= 'sd3289;
        'd1400: dout <= -'sd5234;
        'd1401: dout <= -'sd4560;
        'd1402: dout <= -'sd3096;
        'd1403: dout <= -'sd3722;
        'd1404: dout <= 'sd4479;
        'd1405: dout <= -'sd4070;
        'd1406: dout <= -'sd5203;
        'd1407: dout <= 'sd3109;
        'd1408: dout <= -'sd4736;
        'd1409: dout <= 'sd12;
        'd1410: dout <= 'sd1842;
        'd1411: dout <= -'sd6052;
        'd1412: dout <= -'sd4744;
        'd1413: dout <= -'sd1016;
        'd1414: dout <= 'sd3952;
        'd1415: dout <= -'sd2849;
        'd1416: dout <= 'sd2303;
        'd1417: dout <= -'sd5101;
        'd1418: dout <= 'sd5169;
        'd1419: dout <= -'sd156;
        'd1420: dout <= -'sd2156;
        'd1421: dout <= 'sd3050;
        'd1422: dout <= -'sd374;
        'd1423: dout <= 'sd3029;
        'd1424: dout <= -'sd916;
        'd1425: dout <= -'sd116;
        'd1426: dout <= -'sd3709;
        'd1427: dout <= 'sd718;
        'd1428: dout <= -'sd2627;
        'd1429: dout <= -'sd3328;
        'd1430: dout <= -'sd346;
        'd1431: dout <= 'sd4754;
        'd1432: dout <= -'sd3828;
        'd1433: dout <= 'sd873;
        'd1434: dout <= -'sd1181;
        'd1435: dout <= 'sd103;
        'd1436: dout <= 'sd2;
        'd1437: dout <= -'sd4345;
        'd1438: dout <= 'sd5963;
        'd1439: dout <= -'sd1450;
        'd1440: dout <= -'sd1039;
        'd1441: dout <= -'sd628;
        'd1442: dout <= -'sd747;
        'd1443: dout <= 'sd1382;
        'd1444: dout <= 'sd1257;
        'd1445: dout <= 'sd2666;
        'd1446: dout <= -'sd4998;
        'd1447: dout <= -'sd4389;
        'd1448: dout <= -'sd2906;
        'd1449: dout <= -'sd3977;
        'd1450: dout <= -'sd1254;
        'd1451: dout <= -'sd4799;
        'd1452: dout <= -'sd3018;
        'd1453: dout <= -'sd3;
        'd1454: dout <= 'sd1462;
        'd1455: dout <= -'sd5613;
        'd1456: dout <= -'sd5507;
        'd1457: dout <= 'sd3695;
        'd1458: dout <= 'sd850;
        'd1459: dout <= 'sd1524;
        'd1460: dout <= 'sd3739;
        'd1461: dout <= -'sd3387;
        'd1462: dout <= 'sd4779;
        'd1463: dout <= 'sd1019;
        'd1464: dout <= -'sd1522;
        'd1465: dout <= -'sd5966;
        'd1466: dout <= -'sd5940;
        'd1467: dout <= -'sd4103;
        'd1468: dout <= -'sd5671;
        'd1469: dout <= 'sd5272;
        'd1470: dout <= -'sd1108;
        'd1471: dout <= 'sd4572;
        'd1472: dout <= 'sd4946;
        'd1473: dout <= -'sd2179;
        'd1474: dout <= 'sd4761;
        'd1475: dout <= -'sd5678;
        'd1476: dout <= -'sd476;
        'd1477: dout <= -'sd4468;
        'd1478: dout <= 'sd5003;
        'd1479: dout <= -'sd4932;
        'd1480: dout <= -'sd3348;
        'd1481: dout <= 'sd4986;
        'd1482: dout <= 'sd2349;
        'd1483: dout <= -'sd3587;
        'd1484: dout <= 'sd808;
        'd1485: dout <= 'sd3528;
        'd1486: dout <= -'sd3931;
        'd1487: dout <= -'sd2719;
        'd1488: dout <= -'sd5446;
        'd1489: dout <= -'sd3455;
        'd1490: dout <= 'sd7;
        'd1491: dout <= -'sd2250;
        'd1492: dout <= 'sd4262;
        'd1493: dout <= -'sd2732;
        'd1494: dout <= -'sd1673;
        'd1495: dout <= 'sd859;
        'd1496: dout <= -'sd4852;
        'd1497: dout <= -'sd5095;
        'd1498: dout <= 'sd6107;
        'd1499: dout <= -'sd4375;
        'd1500: dout <= 'sd6043;
        'd1501: dout <= -'sd2420;
        'd1502: dout <= -'sd2800;
        'd1503: dout <= 'sd739;
        'd1504: dout <= 'sd1070;
        'd1505: dout <= -'sd851;
        'd1506: dout <= -'sd320;
        'd1507: dout <= -'sd4463;
        'd1508: dout <= 'sd1476;
        'd1509: dout <= 'sd3937;
        'd1510: dout <= -'sd5956;
        'd1511: dout <= -'sd73;
        'd1512: dout <= -'sd5112;
        'd1513: dout <= -'sd356;
        'd1514: dout <= -'sd5800;
        'd1515: dout <= -'sd5221;
        'd1516: dout <= 'sd3595;
        'd1517: dout <= 'sd71;
        'd1518: dout <= -'sd6044;
        'd1519: dout <= 'sd2214;
        'd1520: dout <= 'sd5712;
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

module hq3_rom (
  input                    clk,
  input                    rst,
  input             [10:0] addr,
  output reg signed [13:0] dout
) ;

  always @ (posedge clk) begin
    if(rst) begin
      dout <= 'sd0;
    end else begin
      case(addr)
        'd0: dout <= -'sd6450;
        'd1: dout <= 'sd167;
        'd2: dout <= 'sd5292;
        'd3: dout <= 'sd6402;
        'd4: dout <= 'sd600;
        'd5: dout <= -'sd788;
        'd6: dout <= -'sd1668;
        'd7: dout <= -'sd7600;
        'd8: dout <= -'sd6471;
        'd9: dout <= -'sd4064;
        'd10: dout <= 'sd3984;
        'd11: dout <= 'sd5148;
        'd12: dout <= 'sd3688;
        'd13: dout <= -'sd3133;
        'd14: dout <= -'sd3070;
        'd15: dout <= -'sd2773;
        'd16: dout <= 'sd4173;
        'd17: dout <= -'sd6643;
        'd18: dout <= 'sd3531;
        'd19: dout <= -'sd4352;
        'd20: dout <= -'sd1484;
        'd21: dout <= 'sd4382;
        'd22: dout <= 'sd2264;
        'd23: dout <= 'sd2868;
        'd24: dout <= 'sd5210;
        'd25: dout <= 'sd1125;
        'd26: dout <= -'sd3704;
        'd27: dout <= 'sd7068;
        'd28: dout <= 'sd3036;
        'd29: dout <= -'sd4509;
        'd30: dout <= -'sd3775;
        'd31: dout <= 'sd1285;
        'd32: dout <= -'sd6834;
        'd33: dout <= -'sd6831;
        'd34: dout <= 'sd5264;
        'd35: dout <= 'sd1254;
        'd36: dout <= -'sd2759;
        'd37: dout <= -'sd7343;
        'd38: dout <= 'sd3726;
        'd39: dout <= -'sd3770;
        'd40: dout <= -'sd3682;
        'd41: dout <= 'sd681;
        'd42: dout <= 'sd3837;
        'd43: dout <= -'sd381;
        'd44: dout <= 'sd5724;
        'd45: dout <= 'sd5852;
        'd46: dout <= 'sd7399;
        'd47: dout <= -'sd7326;
        'd48: dout <= 'sd590;
        'd49: dout <= -'sd7313;
        'd50: dout <= 'sd6225;
        'd51: dout <= 'sd2110;
        'd52: dout <= 'sd679;
        'd53: dout <= -'sd4861;
        'd54: dout <= -'sd1121;
        'd55: dout <= -'sd4865;
        'd56: dout <= 'sd300;
        'd57: dout <= -'sd2264;
        'd58: dout <= 'sd2392;
        'd59: dout <= -'sd1998;
        'd60: dout <= 'sd6020;
        'd61: dout <= -'sd850;
        'd62: dout <= 'sd1034;
        'd63: dout <= 'sd75;
        'd64: dout <= 'sd2256;
        'd65: dout <= -'sd277;
        'd66: dout <= -'sd3838;
        'd67: dout <= -'sd332;
        'd68: dout <= 'sd4903;
        'd69: dout <= -'sd2353;
        'd70: dout <= 'sd5597;
        'd71: dout <= 'sd4436;
        'd72: dout <= -'sd4678;
        'd73: dout <= -'sd4758;
        'd74: dout <= 'sd3007;
        'd75: dout <= -'sd4114;
        'd76: dout <= -'sd730;
        'd77: dout <= 'sd5513;
        'd78: dout <= 'sd1901;
        'd79: dout <= 'sd2332;
        'd80: dout <= -'sd6040;
        'd81: dout <= 'sd1299;
        'd82: dout <= 'sd6236;
        'd83: dout <= -'sd993;
        'd84: dout <= 'sd6555;
        'd85: dout <= -'sd1473;
        'd86: dout <= -'sd868;
        'd87: dout <= 'sd4096;
        'd88: dout <= 'sd191;
        'd89: dout <= 'sd4277;
        'd90: dout <= 'sd2699;
        'd91: dout <= -'sd1728;
        'd92: dout <= 'sd6876;
        'd93: dout <= 'sd310;
        'd94: dout <= -'sd5631;
        'd95: dout <= 'sd1102;
        'd96: dout <= -'sd7120;
        'd97: dout <= -'sd456;
        'd98: dout <= 'sd3425;
        'd99: dout <= 'sd6208;
        'd100: dout <= -'sd5849;
        'd101: dout <= 'sd834;
        'd102: dout <= 'sd1456;
        'd103: dout <= 'sd7184;
        'd104: dout <= 'sd5578;
        'd105: dout <= 'sd6963;
        'd106: dout <= -'sd624;
        'd107: dout <= -'sd4636;
        'd108: dout <= 'sd5252;
        'd109: dout <= 'sd1124;
        'd110: dout <= -'sd2918;
        'd111: dout <= -'sd1485;
        'd112: dout <= -'sd121;
        'd113: dout <= 'sd1965;
        'd114: dout <= 'sd5656;
        'd115: dout <= -'sd7388;
        'd116: dout <= 'sd301;
        'd117: dout <= -'sd1480;
        'd118: dout <= 'sd1318;
        'd119: dout <= -'sd576;
        'd120: dout <= -'sd4624;
        'd121: dout <= -'sd7315;
        'd122: dout <= 'sd2709;
        'd123: dout <= -'sd617;
        'd124: dout <= -'sd3790;
        'd125: dout <= 'sd2635;
        'd126: dout <= 'sd6682;
        'd127: dout <= -'sd4468;
        'd128: dout <= -'sd4012;
        'd129: dout <= -'sd2865;
        'd130: dout <= 'sd3087;
        'd131: dout <= -'sd3284;
        'd132: dout <= 'sd3121;
        'd133: dout <= -'sd2455;
        'd134: dout <= 'sd4149;
        'd135: dout <= -'sd417;
        'd136: dout <= 'sd3397;
        'd137: dout <= 'sd1976;
        'd138: dout <= -'sd7129;
        'd139: dout <= -'sd485;
        'd140: dout <= -'sd522;
        'd141: dout <= -'sd983;
        'd142: dout <= -'sd5360;
        'd143: dout <= 'sd4915;
        'd144: dout <= 'sd4400;
        'd145: dout <= -'sd5141;
        'd146: dout <= 'sd3254;
        'd147: dout <= 'sd636;
        'd148: dout <= 'sd877;
        'd149: dout <= -'sd2004;
        'd150: dout <= -'sd2354;
        'd151: dout <= -'sd4290;
        'd152: dout <= 'sd5686;
        'd153: dout <= -'sd1555;
        'd154: dout <= -'sd6675;
        'd155: dout <= -'sd4040;
        'd156: dout <= -'sd727;
        'd157: dout <= 'sd5244;
        'd158: dout <= -'sd5500;
        'd159: dout <= 'sd7014;
        'd160: dout <= -'sd6561;
        'd161: dout <= 'sd378;
        'd162: dout <= 'sd709;
        'd163: dout <= -'sd7419;
        'd164: dout <= -'sd405;
        'd165: dout <= 'sd4814;
        'd166: dout <= 'sd5433;
        'd167: dout <= 'sd501;
        'd168: dout <= 'sd4611;
        'd169: dout <= -'sd1532;
        'd170: dout <= -'sd6100;
        'd171: dout <= -'sd1496;
        'd172: dout <= 'sd7452;
        'd173: dout <= -'sd4790;
        'd174: dout <= -'sd3916;
        'd175: dout <= 'sd6657;
        'd176: dout <= 'sd4552;
        'd177: dout <= -'sd6744;
        'd178: dout <= 'sd5836;
        'd179: dout <= 'sd2553;
        'd180: dout <= -'sd3758;
        'd181: dout <= 'sd202;
        'd182: dout <= -'sd1492;
        'd183: dout <= 'sd6323;
        'd184: dout <= 'sd7433;
        'd185: dout <= -'sd3844;
        'd186: dout <= 'sd1979;
        'd187: dout <= 'sd3189;
        'd188: dout <= -'sd1555;
        'd189: dout <= 'sd4873;
        'd190: dout <= -'sd436;
        'd191: dout <= 'sd3759;
        'd192: dout <= 'sd6747;
        'd193: dout <= -'sd2287;
        'd194: dout <= 'sd4843;
        'd195: dout <= -'sd6379;
        'd196: dout <= 'sd472;
        'd197: dout <= 'sd4231;
        'd198: dout <= -'sd7392;
        'd199: dout <= 'sd5638;
        'd200: dout <= 'sd2120;
        'd201: dout <= -'sd1668;
        'd202: dout <= -'sd3544;
        'd203: dout <= 'sd2001;
        'd204: dout <= 'sd1959;
        'd205: dout <= -'sd3204;
        'd206: dout <= 'sd326;
        'd207: dout <= -'sd5263;
        'd208: dout <= -'sd5735;
        'd209: dout <= -'sd3318;
        'd210: dout <= 'sd245;
        'd211: dout <= 'sd6837;
        'd212: dout <= 'sd4250;
        'd213: dout <= 'sd365;
        'd214: dout <= 'sd3113;
        'd215: dout <= 'sd3377;
        'd216: dout <= 'sd1154;
        'd217: dout <= -'sd7620;
        'd218: dout <= -'sd4139;
        'd219: dout <= 'sd1303;
        'd220: dout <= 'sd6204;
        'd221: dout <= 'sd5164;
        'd222: dout <= -'sd5417;
        'd223: dout <= 'sd7157;
        'd224: dout <= -'sd1367;
        'd225: dout <= 'sd3964;
        'd226: dout <= 'sd6576;
        'd227: dout <= -'sd2381;
        'd228: dout <= -'sd3678;
        'd229: dout <= 'sd4663;
        'd230: dout <= -'sd3826;
        'd231: dout <= 'sd3283;
        'd232: dout <= -'sd7518;
        'd233: dout <= 'sd2479;
        'd234: dout <= 'sd6321;
        'd235: dout <= 'sd5227;
        'd236: dout <= 'sd5804;
        'd237: dout <= 'sd6775;
        'd238: dout <= 'sd6384;
        'd239: dout <= -'sd6959;
        'd240: dout <= 'sd4327;
        'd241: dout <= -'sd2349;
        'd242: dout <= -'sd565;
        'd243: dout <= 'sd125;
        'd244: dout <= -'sd256;
        'd245: dout <= 'sd5237;
        'd246: dout <= 'sd6515;
        'd247: dout <= 'sd5144;
        'd248: dout <= -'sd6365;
        'd249: dout <= -'sd4148;
        'd250: dout <= -'sd2967;
        'd251: dout <= 'sd4612;
        'd252: dout <= 'sd400;
        'd253: dout <= 'sd4225;
        'd254: dout <= 'sd117;
        'd255: dout <= 'sd1303;
        'd256: dout <= -'sd4834;
        'd257: dout <= 'sd806;
        'd258: dout <= -'sd4816;
        'd259: dout <= -'sd2622;
        'd260: dout <= 'sd1296;
        'd261: dout <= -'sd448;
        'd262: dout <= 'sd6349;
        'd263: dout <= -'sd1827;
        'd264: dout <= -'sd5113;
        'd265: dout <= 'sd7273;
        'd266: dout <= -'sd1773;
        'd267: dout <= -'sd2399;
        'd268: dout <= 'sd1578;
        'd269: dout <= 'sd3748;
        'd270: dout <= -'sd2797;
        'd271: dout <= 'sd585;
        'd272: dout <= -'sd3019;
        'd273: dout <= 'sd1318;
        'd274: dout <= -'sd1296;
        'd275: dout <= -'sd5034;
        'd276: dout <= 'sd279;
        'd277: dout <= -'sd1682;
        'd278: dout <= 'sd1975;
        'd279: dout <= 'sd1034;
        'd280: dout <= -'sd6909;
        'd281: dout <= 'sd110;
        'd282: dout <= -'sd7084;
        'd283: dout <= -'sd2422;
        'd284: dout <= 'sd7018;
        'd285: dout <= -'sd7460;
        'd286: dout <= 'sd7355;
        'd287: dout <= 'sd3008;
        'd288: dout <= -'sd3393;
        'd289: dout <= 'sd18;
        'd290: dout <= -'sd1156;
        'd291: dout <= 'sd1631;
        'd292: dout <= 'sd5990;
        'd293: dout <= 'sd2150;
        'd294: dout <= -'sd6002;
        'd295: dout <= 'sd3884;
        'd296: dout <= 'sd7637;
        'd297: dout <= -'sd605;
        'd298: dout <= 'sd7202;
        'd299: dout <= -'sd2355;
        'd300: dout <= 'sd889;
        'd301: dout <= -'sd242;
        'd302: dout <= 'sd2975;
        'd303: dout <= 'sd3164;
        'd304: dout <= -'sd4975;
        'd305: dout <= -'sd1973;
        'd306: dout <= -'sd6769;
        'd307: dout <= -'sd6524;
        'd308: dout <= -'sd5950;
        'd309: dout <= 'sd5418;
        'd310: dout <= 'sd5577;
        'd311: dout <= -'sd3546;
        'd312: dout <= -'sd5311;
        'd313: dout <= -'sd7593;
        'd314: dout <= 'sd6379;
        'd315: dout <= 'sd2294;
        'd316: dout <= -'sd2687;
        'd317: dout <= -'sd4486;
        'd318: dout <= 'sd731;
        'd319: dout <= -'sd2159;
        'd320: dout <= -'sd947;
        'd321: dout <= -'sd6732;
        'd322: dout <= -'sd833;
        'd323: dout <= -'sd2789;
        'd324: dout <= -'sd989;
        'd325: dout <= -'sd1756;
        'd326: dout <= -'sd3646;
        'd327: dout <= -'sd4207;
        'd328: dout <= -'sd6629;
        'd329: dout <= -'sd7513;
        'd330: dout <= 'sd5919;
        'd331: dout <= 'sd3670;
        'd332: dout <= 'sd1496;
        'd333: dout <= -'sd6707;
        'd334: dout <= 'sd6684;
        'd335: dout <= 'sd1337;
        'd336: dout <= -'sd6279;
        'd337: dout <= 'sd2380;
        'd338: dout <= 'sd2525;
        'd339: dout <= 'sd3696;
        'd340: dout <= 'sd3249;
        'd341: dout <= -'sd7009;
        'd342: dout <= -'sd4852;
        'd343: dout <= -'sd1765;
        'd344: dout <= -'sd2112;
        'd345: dout <= -'sd4361;
        'd346: dout <= 'sd140;
        'd347: dout <= -'sd634;
        'd348: dout <= -'sd4921;
        'd349: dout <= 'sd6388;
        'd350: dout <= -'sd846;
        'd351: dout <= 'sd5931;
        'd352: dout <= -'sd1564;
        'd353: dout <= -'sd7264;
        'd354: dout <= -'sd4464;
        'd355: dout <= -'sd475;
        'd356: dout <= 'sd5310;
        'd357: dout <= -'sd2970;
        'd358: dout <= -'sd4373;
        'd359: dout <= -'sd4522;
        'd360: dout <= -'sd4511;
        'd361: dout <= 'sd5421;
        'd362: dout <= -'sd114;
        'd363: dout <= -'sd1154;
        'd364: dout <= 'sd7370;
        'd365: dout <= -'sd1052;
        'd366: dout <= 'sd7166;
        'd367: dout <= -'sd5176;
        'd368: dout <= -'sd4891;
        'd369: dout <= 'sd4984;
        'd370: dout <= 'sd4608;
        'd371: dout <= -'sd906;
        'd372: dout <= 'sd7090;
        'd373: dout <= 'sd5836;
        'd374: dout <= 'sd2917;
        'd375: dout <= 'sd4688;
        'd376: dout <= -'sd178;
        'd377: dout <= -'sd122;
        'd378: dout <= 'sd6985;
        'd379: dout <= -'sd2090;
        'd380: dout <= -'sd5036;
        'd381: dout <= -'sd4183;
        'd382: dout <= -'sd1967;
        'd383: dout <= 'sd7263;
        'd384: dout <= -'sd2481;
        'd385: dout <= -'sd3428;
        'd386: dout <= 'sd5038;
        'd387: dout <= -'sd3906;
        'd388: dout <= -'sd5714;
        'd389: dout <= 'sd2062;
        'd390: dout <= 'sd4545;
        'd391: dout <= -'sd4775;
        'd392: dout <= 'sd1841;
        'd393: dout <= -'sd3763;
        'd394: dout <= -'sd313;
        'd395: dout <= 'sd437;
        'd396: dout <= -'sd2459;
        'd397: dout <= 'sd1971;
        'd398: dout <= 'sd5997;
        'd399: dout <= 'sd7522;
        'd400: dout <= -'sd3036;
        'd401: dout <= 'sd1399;
        'd402: dout <= 'sd5826;
        'd403: dout <= 'sd4159;
        'd404: dout <= 'sd1672;
        'd405: dout <= 'sd6250;
        'd406: dout <= -'sd247;
        'd407: dout <= 'sd1465;
        'd408: dout <= 'sd3325;
        'd409: dout <= -'sd1080;
        'd410: dout <= 'sd1548;
        'd411: dout <= 'sd3483;
        'd412: dout <= -'sd358;
        'd413: dout <= 'sd2420;
        'd414: dout <= -'sd3556;
        'd415: dout <= -'sd5244;
        'd416: dout <= -'sd4701;
        'd417: dout <= -'sd7508;
        'd418: dout <= 'sd2837;
        'd419: dout <= 'sd1225;
        'd420: dout <= -'sd3916;
        'd421: dout <= -'sd6978;
        'd422: dout <= -'sd5365;
        'd423: dout <= -'sd3281;
        'd424: dout <= -'sd6706;
        'd425: dout <= 'sd2490;
        'd426: dout <= -'sd6219;
        'd427: dout <= -'sd6389;
        'd428: dout <= 'sd6083;
        'd429: dout <= -'sd2161;
        'd430: dout <= -'sd75;
        'd431: dout <= -'sd2458;
        'd432: dout <= -'sd1539;
        'd433: dout <= -'sd5450;
        'd434: dout <= 'sd3540;
        'd435: dout <= 'sd4449;
        'd436: dout <= 'sd1516;
        'd437: dout <= 'sd7050;
        'd438: dout <= 'sd1238;
        'd439: dout <= 'sd6461;
        'd440: dout <= 'sd2388;
        'd441: dout <= -'sd3715;
        'd442: dout <= 'sd5386;
        'd443: dout <= 'sd4304;
        'd444: dout <= -'sd4394;
        'd445: dout <= -'sd3776;
        'd446: dout <= -'sd2992;
        'd447: dout <= 'sd744;
        'd448: dout <= 'sd5616;
        'd449: dout <= -'sd4822;
        'd450: dout <= 'sd637;
        'd451: dout <= -'sd5693;
        'd452: dout <= 'sd820;
        'd453: dout <= -'sd7277;
        'd454: dout <= -'sd4303;
        'd455: dout <= -'sd2225;
        'd456: dout <= 'sd1815;
        'd457: dout <= 'sd6643;
        'd458: dout <= -'sd1733;
        'd459: dout <= 'sd6809;
        'd460: dout <= -'sd2557;
        'd461: dout <= 'sd6837;
        'd462: dout <= 'sd1315;
        'd463: dout <= 'sd4434;
        'd464: dout <= 'sd4590;
        'd465: dout <= 'sd63;
        'd466: dout <= -'sd2849;
        'd467: dout <= 'sd2822;
        'd468: dout <= 'sd970;
        'd469: dout <= 'sd3509;
        'd470: dout <= -'sd6537;
        'd471: dout <= 'sd3687;
        'd472: dout <= 'sd5784;
        'd473: dout <= -'sd1931;
        'd474: dout <= -'sd2408;
        'd475: dout <= 'sd4050;
        'd476: dout <= 'sd3091;
        'd477: dout <= 'sd1976;
        'd478: dout <= -'sd1511;
        'd479: dout <= 'sd816;
        'd480: dout <= -'sd2208;
        'd481: dout <= -'sd6218;
        'd482: dout <= 'sd6285;
        'd483: dout <= -'sd3769;
        'd484: dout <= 'sd4586;
        'd485: dout <= 'sd6092;
        'd486: dout <= 'sd6468;
        'd487: dout <= -'sd5068;
        'd488: dout <= 'sd1371;
        'd489: dout <= -'sd5021;
        'd490: dout <= 'sd2229;
        'd491: dout <= -'sd4867;
        'd492: dout <= 'sd3212;
        'd493: dout <= 'sd1526;
        'd494: dout <= -'sd3539;
        'd495: dout <= -'sd3072;
        'd496: dout <= -'sd1528;
        'd497: dout <= 'sd7501;
        'd498: dout <= 'sd2771;
        'd499: dout <= 'sd2122;
        'd500: dout <= -'sd7633;
        'd501: dout <= 'sd892;
        'd502: dout <= -'sd1140;
        'd503: dout <= 'sd5319;
        'd504: dout <= -'sd1666;
        'd505: dout <= -'sd477;
        'd506: dout <= -'sd3011;
        'd507: dout <= -'sd939;
        'd508: dout <= 'sd1305;
        'd509: dout <= -'sd4623;
        'd510: dout <= 'sd7404;
        'd511: dout <= -'sd5737;
        'd512: dout <= 'sd951;
        'd513: dout <= 'sd6037;
        'd514: dout <= 'sd5910;
        'd515: dout <= -'sd924;
        'd516: dout <= 'sd2451;
        'd517: dout <= -'sd5295;
        'd518: dout <= -'sd3492;
        'd519: dout <= -'sd2062;
        'd520: dout <= -'sd6268;
        'd521: dout <= -'sd3306;
        'd522: dout <= -'sd6388;
        'd523: dout <= 'sd2311;
        'd524: dout <= -'sd1639;
        'd525: dout <= -'sd4569;
        'd526: dout <= 'sd890;
        'd527: dout <= -'sd6790;
        'd528: dout <= 'sd834;
        'd529: dout <= -'sd1551;
        'd530: dout <= -'sd7672;
        'd531: dout <= -'sd6625;
        'd532: dout <= 'sd7185;
        'd533: dout <= 'sd3343;
        'd534: dout <= -'sd4248;
        'd535: dout <= -'sd2649;
        'd536: dout <= 'sd7485;
        'd537: dout <= 'sd2869;
        'd538: dout <= 'sd7283;
        'd539: dout <= -'sd4151;
        'd540: dout <= -'sd2147;
        'd541: dout <= 'sd5948;
        'd542: dout <= 'sd3484;
        'd543: dout <= 'sd5895;
        'd544: dout <= -'sd7287;
        'd545: dout <= -'sd6933;
        'd546: dout <= -'sd820;
        'd547: dout <= -'sd22;
        'd548: dout <= -'sd617;
        'd549: dout <= 'sd5261;
        'd550: dout <= 'sd1868;
        'd551: dout <= 'sd2796;
        'd552: dout <= 'sd6570;
        'd553: dout <= -'sd4301;
        'd554: dout <= -'sd6292;
        'd555: dout <= 'sd2644;
        'd556: dout <= 'sd5751;
        'd557: dout <= 'sd2676;
        'd558: dout <= -'sd3905;
        'd559: dout <= -'sd1926;
        'd560: dout <= 'sd1075;
        'd561: dout <= -'sd1528;
        'd562: dout <= 'sd1703;
        'd563: dout <= -'sd2077;
        'd564: dout <= -'sd2753;
        'd565: dout <= -'sd6551;
        'd566: dout <= 'sd2396;
        'd567: dout <= -'sd6241;
        'd568: dout <= -'sd6618;
        'd569: dout <= 'sd3812;
        'd570: dout <= 'sd6490;
        'd571: dout <= -'sd6570;
        'd572: dout <= -'sd6223;
        'd573: dout <= 'sd5175;
        'd574: dout <= -'sd6254;
        'd575: dout <= -'sd3511;
        'd576: dout <= 'sd3520;
        'd577: dout <= 'sd5303;
        'd578: dout <= 'sd4505;
        'd579: dout <= -'sd329;
        'd580: dout <= -'sd7388;
        'd581: dout <= -'sd5013;
        'd582: dout <= -'sd3952;
        'd583: dout <= -'sd4385;
        'd584: dout <= -'sd1962;
        'd585: dout <= -'sd6870;
        'd586: dout <= 'sd2217;
        'd587: dout <= 'sd1613;
        'd588: dout <= -'sd7571;
        'd589: dout <= 'sd3372;
        'd590: dout <= -'sd5541;
        'd591: dout <= 'sd2044;
        'd592: dout <= 'sd7674;
        'd593: dout <= 'sd3871;
        'd594: dout <= 'sd4584;
        'd595: dout <= -'sd4763;
        'd596: dout <= -'sd1825;
        'd597: dout <= -'sd7127;
        'd598: dout <= -'sd449;
        'd599: dout <= -'sd380;
        'd600: dout <= -'sd337;
        'd601: dout <= 'sd4075;
        'd602: dout <= -'sd1102;
        'd603: dout <= -'sd3487;
        'd604: dout <= -'sd47;
        'd605: dout <= -'sd2243;
        'd606: dout <= -'sd996;
        'd607: dout <= -'sd5297;
        'd608: dout <= -'sd3020;
        'd609: dout <= 'sd5620;
        'd610: dout <= -'sd7243;
        'd611: dout <= 'sd432;
        'd612: dout <= 'sd4633;
        'd613: dout <= -'sd1580;
        'd614: dout <= 'sd3736;
        'd615: dout <= 'sd630;
        'd616: dout <= -'sd5464;
        'd617: dout <= -'sd6628;
        'd618: dout <= 'sd187;
        'd619: dout <= -'sd5908;
        'd620: dout <= 'sd1519;
        'd621: dout <= -'sd7234;
        'd622: dout <= -'sd3372;
        'd623: dout <= 'sd2217;
        'd624: dout <= 'sd3035;
        'd625: dout <= 'sd5456;
        'd626: dout <= -'sd6261;
        'd627: dout <= -'sd1455;
        'd628: dout <= -'sd2448;
        'd629: dout <= -'sd875;
        'd630: dout <= 'sd5906;
        'd631: dout <= 'sd6262;
        'd632: dout <= -'sd6764;
        'd633: dout <= -'sd3659;
        'd634: dout <= 'sd1923;
        'd635: dout <= -'sd3215;
        'd636: dout <= 'sd6255;
        'd637: dout <= -'sd2418;
        'd638: dout <= 'sd6276;
        'd639: dout <= 'sd5328;
        'd640: dout <= -'sd7251;
        'd641: dout <= 'sd4187;
        'd642: dout <= -'sd1027;
        'd643: dout <= -'sd3709;
        'd644: dout <= -'sd4183;
        'd645: dout <= 'sd5379;
        'd646: dout <= -'sd6232;
        'd647: dout <= 'sd3794;
        'd648: dout <= 'sd5316;
        'd649: dout <= 'sd6901;
        'd650: dout <= -'sd5350;
        'd651: dout <= -'sd2409;
        'd652: dout <= 'sd1658;
        'd653: dout <= -'sd4583;
        'd654: dout <= 'sd1237;
        'd655: dout <= -'sd6010;
        'd656: dout <= -'sd2408;
        'd657: dout <= 'sd3088;
        'd658: dout <= -'sd6320;
        'd659: dout <= -'sd5288;
        'd660: dout <= -'sd7495;
        'd661: dout <= 'sd5028;
        'd662: dout <= 'sd7571;
        'd663: dout <= 'sd4125;
        'd664: dout <= 'sd7397;
        'd665: dout <= 'sd325;
        'd666: dout <= -'sd2316;
        'd667: dout <= 'sd3932;
        'd668: dout <= 'sd431;
        'd669: dout <= 'sd2256;
        'd670: dout <= -'sd3206;
        'd671: dout <= 'sd682;
        'd672: dout <= -'sd6176;
        'd673: dout <= -'sd5343;
        'd674: dout <= 'sd3915;
        'd675: dout <= -'sd2078;
        'd676: dout <= 'sd1754;
        'd677: dout <= -'sd6337;
        'd678: dout <= -'sd6103;
        'd679: dout <= -'sd7487;
        'd680: dout <= -'sd2823;
        'd681: dout <= -'sd1933;
        'd682: dout <= -'sd2485;
        'd683: dout <= 'sd5967;
        'd684: dout <= -'sd2050;
        'd685: dout <= 'sd1411;
        'd686: dout <= -'sd2492;
        'd687: dout <= -'sd3486;
        'd688: dout <= -'sd5653;
        'd689: dout <= -'sd3423;
        'd690: dout <= 'sd4074;
        'd691: dout <= 'sd3359;
        'd692: dout <= 'sd3588;
        'd693: dout <= -'sd69;
        'd694: dout <= 'sd6223;
        'd695: dout <= 'sd1977;
        'd696: dout <= -'sd6396;
        'd697: dout <= -'sd402;
        'd698: dout <= -'sd1729;
        'd699: dout <= 'sd4336;
        'd700: dout <= -'sd4540;
        'd701: dout <= -'sd6022;
        'd702: dout <= -'sd1827;
        'd703: dout <= 'sd4959;
        'd704: dout <= -'sd6743;
        'd705: dout <= -'sd5554;
        'd706: dout <= -'sd4639;
        'd707: dout <= 'sd4641;
        'd708: dout <= -'sd4590;
        'd709: dout <= -'sd3656;
        'd710: dout <= -'sd1146;
        'd711: dout <= -'sd3940;
        'd712: dout <= 'sd2846;
        'd713: dout <= 'sd4960;
        'd714: dout <= 'sd1717;
        'd715: dout <= 'sd3355;
        'd716: dout <= 'sd5770;
        'd717: dout <= 'sd7098;
        'd718: dout <= -'sd664;
        'd719: dout <= -'sd7102;
        'd720: dout <= -'sd2438;
        'd721: dout <= -'sd2504;
        'd722: dout <= -'sd1258;
        'd723: dout <= -'sd2771;
        'd724: dout <= 'sd3279;
        'd725: dout <= -'sd6742;
        'd726: dout <= -'sd2554;
        'd727: dout <= 'sd214;
        'd728: dout <= -'sd3250;
        'd729: dout <= -'sd5382;
        'd730: dout <= -'sd7525;
        'd731: dout <= -'sd6270;
        'd732: dout <= 'sd5243;
        'd733: dout <= -'sd4473;
        'd734: dout <= -'sd3310;
        'd735: dout <= 'sd3770;
        'd736: dout <= 'sd2775;
        'd737: dout <= -'sd1435;
        'd738: dout <= 'sd3862;
        'd739: dout <= -'sd1228;
        'd740: dout <= -'sd7085;
        'd741: dout <= -'sd3043;
        'd742: dout <= 'sd4209;
        'd743: dout <= 'sd830;
        'd744: dout <= -'sd4832;
        'd745: dout <= -'sd3314;
        'd746: dout <= -'sd1440;
        'd747: dout <= 'sd5938;
        'd748: dout <= 'sd5427;
        'd749: dout <= -'sd6576;
        'd750: dout <= -'sd408;
        'd751: dout <= 'sd3001;
        'd752: dout <= -'sd4445;
        'd753: dout <= 'sd2173;
        'd754: dout <= -'sd6263;
        'd755: dout <= -'sd2866;
        'd756: dout <= -'sd3187;
        'd757: dout <= 'sd851;
        'd758: dout <= 'sd2392;
        'd759: dout <= -'sd1051;
        'd760: dout <= -'sd6286;
        'd761: dout <= -'sd2313;
        'd762: dout <= -'sd1619;
        'd763: dout <= -'sd305;
        'd764: dout <= 'sd1503;
        'd765: dout <= -'sd7296;
        'd766: dout <= -'sd1705;
        'd767: dout <= 'sd438;
        'd768: dout <= 'sd3384;
        'd769: dout <= -'sd7601;
        'd770: dout <= -'sd2226;
        'd771: dout <= 'sd3239;
        'd772: dout <= -'sd2317;
        'd773: dout <= 'sd6771;
        'd774: dout <= 'sd2269;
        'd775: dout <= 'sd2291;
        'd776: dout <= -'sd4193;
        'd777: dout <= -'sd5014;
        'd778: dout <= 'sd3475;
        'd779: dout <= -'sd2051;
        'd780: dout <= -'sd2538;
        'd781: dout <= 'sd1173;
        'd782: dout <= 'sd3504;
        'd783: dout <= -'sd25;
        'd784: dout <= 'sd6589;
        'd785: dout <= 'sd4332;
        'd786: dout <= 'sd104;
        'd787: dout <= -'sd5961;
        'd788: dout <= 'sd1024;
        'd789: dout <= 'sd5242;
        'd790: dout <= 'sd5539;
        'd791: dout <= 'sd6964;
        'd792: dout <= -'sd5813;
        'd793: dout <= -'sd4331;
        'd794: dout <= -'sd3159;
        'd795: dout <= 'sd4652;
        'd796: dout <= 'sd7542;
        'd797: dout <= -'sd3075;
        'd798: dout <= -'sd2064;
        'd799: dout <= -'sd196;
        'd800: dout <= 'sd5660;
        'd801: dout <= 'sd5963;
        'd802: dout <= 'sd384;
        'd803: dout <= -'sd449;
        'd804: dout <= 'sd969;
        'd805: dout <= 'sd6219;
        'd806: dout <= -'sd686;
        'd807: dout <= 'sd4088;
        'd808: dout <= -'sd515;
        'd809: dout <= -'sd6371;
        'd810: dout <= -'sd7339;
        'd811: dout <= 'sd240;
        'd812: dout <= 'sd6707;
        'd813: dout <= 'sd88;
        'd814: dout <= -'sd2337;
        'd815: dout <= -'sd1614;
        'd816: dout <= 'sd7130;
        'd817: dout <= 'sd6479;
        'd818: dout <= 'sd2908;
        'd819: dout <= -'sd269;
        'd820: dout <= -'sd737;
        'd821: dout <= -'sd5044;
        'd822: dout <= -'sd1979;
        'd823: dout <= 'sd5741;
        'd824: dout <= 'sd4526;
        'd825: dout <= -'sd4516;
        'd826: dout <= -'sd6445;
        'd827: dout <= 'sd2028;
        'd828: dout <= -'sd7585;
        'd829: dout <= 'sd1859;
        'd830: dout <= 'sd4600;
        'd831: dout <= -'sd3752;
        'd832: dout <= -'sd4460;
        'd833: dout <= 'sd5507;
        'd834: dout <= 'sd5306;
        'd835: dout <= -'sd4359;
        'd836: dout <= 'sd2858;
        'd837: dout <= 'sd4022;
        'd838: dout <= 'sd45;
        'd839: dout <= 'sd1557;
        'd840: dout <= 'sd3615;
        'd841: dout <= 'sd4407;
        'd842: dout <= 'sd5634;
        'd843: dout <= -'sd685;
        'd844: dout <= -'sd2617;
        'd845: dout <= -'sd4533;
        'd846: dout <= -'sd4537;
        'd847: dout <= -'sd2974;
        'd848: dout <= 'sd7508;
        'd849: dout <= -'sd7307;
        'd850: dout <= -'sd6487;
        'd851: dout <= 'sd7340;
        'd852: dout <= 'sd1914;
        'd853: dout <= 'sd1751;
        'd854: dout <= -'sd6883;
        'd855: dout <= -'sd5685;
        'd856: dout <= 'sd1021;
        'd857: dout <= -'sd5281;
        'd858: dout <= -'sd38;
        'd859: dout <= 'sd3372;
        'd860: dout <= -'sd3952;
        'd861: dout <= 'sd2329;
        'd862: dout <= 'sd7057;
        'd863: dout <= 'sd4466;
        'd864: dout <= -'sd5362;
        'd865: dout <= 'sd5715;
        'd866: dout <= 'sd841;
        'd867: dout <= 'sd3595;
        'd868: dout <= 'sd768;
        'd869: dout <= -'sd822;
        'd870: dout <= 'sd1958;
        'd871: dout <= -'sd6558;
        'd872: dout <= 'sd4910;
        'd873: dout <= 'sd2477;
        'd874: dout <= 'sd1321;
        'd875: dout <= -'sd907;
        'd876: dout <= -'sd290;
        'd877: dout <= -'sd3017;
        'd878: dout <= 'sd754;
        'd879: dout <= -'sd4409;
        'd880: dout <= 'sd3982;
        'd881: dout <= 'sd3118;
        'd882: dout <= -'sd6863;
        'd883: dout <= -'sd4641;
        'd884: dout <= -'sd3137;
        'd885: dout <= 'sd290;
        'd886: dout <= -'sd2636;
        'd887: dout <= 'sd4607;
        'd888: dout <= -'sd2327;
        'd889: dout <= -'sd3275;
        'd890: dout <= 'sd5564;
        'd891: dout <= -'sd3678;
        'd892: dout <= 'sd893;
        'd893: dout <= -'sd439;
        'd894: dout <= 'sd5407;
        'd895: dout <= -'sd4164;
        'd896: dout <= -'sd2287;
        'd897: dout <= -'sd983;
        'd898: dout <= -'sd3763;
        'd899: dout <= 'sd1528;
        'd900: dout <= -'sd4568;
        'd901: dout <= -'sd5171;
        'd902: dout <= 'sd6929;
        'd903: dout <= 'sd4527;
        'd904: dout <= -'sd2355;
        'd905: dout <= 'sd4286;
        'd906: dout <= 'sd3044;
        'd907: dout <= -'sd1083;
        'd908: dout <= 'sd165;
        'd909: dout <= 'sd3000;
        'd910: dout <= 'sd6151;
        'd911: dout <= -'sd7298;
        'd912: dout <= 'sd4740;
        'd913: dout <= -'sd559;
        'd914: dout <= -'sd2691;
        'd915: dout <= 'sd645;
        'd916: dout <= 'sd1852;
        'd917: dout <= 'sd4352;
        'd918: dout <= -'sd2240;
        'd919: dout <= 'sd4850;
        'd920: dout <= 'sd196;
        'd921: dout <= 'sd4955;
        'd922: dout <= 'sd3787;
        'd923: dout <= -'sd6637;
        'd924: dout <= 'sd2580;
        'd925: dout <= 'sd1108;
        'd926: dout <= -'sd3408;
        'd927: dout <= -'sd3604;
        'd928: dout <= 'sd392;
        'd929: dout <= -'sd4668;
        'd930: dout <= -'sd6500;
        'd931: dout <= -'sd4666;
        'd932: dout <= 'sd3037;
        'd933: dout <= -'sd2332;
        'd934: dout <= -'sd215;
        'd935: dout <= -'sd6911;
        'd936: dout <= -'sd5643;
        'd937: dout <= -'sd4488;
        'd938: dout <= -'sd255;
        'd939: dout <= 'sd5187;
        'd940: dout <= -'sd649;
        'd941: dout <= -'sd2500;
        'd942: dout <= 'sd6613;
        'd943: dout <= -'sd4544;
        'd944: dout <= -'sd3029;
        'd945: dout <= 'sd2944;
        'd946: dout <= -'sd4313;
        'd947: dout <= 'sd5488;
        'd948: dout <= 'sd3482;
        'd949: dout <= -'sd6632;
        'd950: dout <= -'sd4987;
        'd951: dout <= 'sd4559;
        'd952: dout <= 'sd7093;
        'd953: dout <= -'sd5367;
        'd954: dout <= 'sd5970;
        'd955: dout <= 'sd2382;
        'd956: dout <= -'sd3568;
        'd957: dout <= 'sd5469;
        'd958: dout <= -'sd1679;
        'd959: dout <= -'sd5436;
        'd960: dout <= 'sd2544;
        'd961: dout <= -'sd897;
        'd962: dout <= -'sd2813;
        'd963: dout <= 'sd4871;
        'd964: dout <= -'sd178;
        'd965: dout <= -'sd7142;
        'd966: dout <= -'sd1679;
        'd967: dout <= 'sd1415;
        'd968: dout <= 'sd349;
        'd969: dout <= 'sd1486;
        'd970: dout <= -'sd5710;
        'd971: dout <= 'sd4655;
        'd972: dout <= 'sd2900;
        'd973: dout <= -'sd75;
        'd974: dout <= 'sd4589;
        'd975: dout <= 'sd3478;
        'd976: dout <= -'sd5023;
        'd977: dout <= -'sd3021;
        'd978: dout <= 'sd1611;
        'd979: dout <= -'sd5880;
        'd980: dout <= 'sd7187;
        'd981: dout <= 'sd7007;
        'd982: dout <= -'sd526;
        'd983: dout <= 'sd3202;
        'd984: dout <= 'sd730;
        'd985: dout <= -'sd1099;
        'd986: dout <= 'sd771;
        'd987: dout <= -'sd7553;
        'd988: dout <= 'sd6723;
        'd989: dout <= -'sd3992;
        'd990: dout <= -'sd1106;
        'd991: dout <= -'sd3359;
        'd992: dout <= 'sd1056;
        'd993: dout <= 'sd3764;
        'd994: dout <= 'sd6066;
        'd995: dout <= 'sd6667;
        'd996: dout <= -'sd6068;
        'd997: dout <= -'sd7075;
        'd998: dout <= -'sd6211;
        'd999: dout <= 'sd2831;
        'd1000: dout <= 'sd432;
        'd1001: dout <= -'sd2320;
        'd1002: dout <= 'sd3475;
        'd1003: dout <= -'sd5274;
        'd1004: dout <= 'sd7373;
        'd1005: dout <= -'sd5697;
        'd1006: dout <= -'sd1130;
        'd1007: dout <= 'sd6784;
        'd1008: dout <= 'sd2444;
        'd1009: dout <= 'sd4448;
        'd1010: dout <= 'sd5274;
        'd1011: dout <= 'sd630;
        'd1012: dout <= -'sd1146;
        'd1013: dout <= 'sd5282;
        'd1014: dout <= 'sd3046;
        'd1015: dout <= 'sd3935;
        'd1016: dout <= 'sd389;
        'd1017: dout <= -'sd703;
        'd1018: dout <= 'sd2982;
        'd1019: dout <= 'sd6377;
        'd1020: dout <= 'sd2779;
        'd1021: dout <= -'sd7285;
        'd1022: dout <= 'sd4897;
        'd1023: dout <= 'sd90;
        'd1024: dout <= 'sd4093;
        'd1025: dout <= -'sd1158;
        'd1026: dout <= 'sd3301;
        'd1027: dout <= 'sd945;
        'd1028: dout <= 'sd524;
        'd1029: dout <= 'sd6164;
        'd1030: dout <= 'sd6517;
        'd1031: dout <= -'sd6175;
        'd1032: dout <= 'sd1;
        'd1033: dout <= -'sd1520;
        'd1034: dout <= -'sd2040;
        'd1035: dout <= 'sd4836;
        'd1036: dout <= -'sd6021;
        'd1037: dout <= 'sd5446;
        'd1038: dout <= 'sd6483;
        'd1039: dout <= -'sd3807;
        'd1040: dout <= 'sd7357;
        'd1041: dout <= 'sd649;
        'd1042: dout <= -'sd3644;
        'd1043: dout <= -'sd3805;
        'd1044: dout <= -'sd6628;
        'd1045: dout <= 'sd7119;
        'd1046: dout <= -'sd6505;
        'd1047: dout <= 'sd2650;
        'd1048: dout <= 'sd4881;
        'd1049: dout <= 'sd3709;
        'd1050: dout <= 'sd6988;
        'd1051: dout <= -'sd4971;
        'd1052: dout <= 'sd5646;
        'd1053: dout <= -'sd3247;
        'd1054: dout <= 'sd5098;
        'd1055: dout <= 'sd4980;
        'd1056: dout <= -'sd6894;
        'd1057: dout <= 'sd5597;
        'd1058: dout <= -'sd7212;
        'd1059: dout <= -'sd5359;
        'd1060: dout <= -'sd1966;
        'd1061: dout <= 'sd3153;
        'd1062: dout <= 'sd6608;
        'd1063: dout <= 'sd4049;
        'd1064: dout <= -'sd5595;
        'd1065: dout <= 'sd4251;
        'd1066: dout <= 'sd1778;
        'd1067: dout <= -'sd1601;
        'd1068: dout <= 'sd2070;
        'd1069: dout <= 'sd6244;
        'd1070: dout <= 'sd1005;
        'd1071: dout <= 'sd637;
        'd1072: dout <= -'sd7420;
        'd1073: dout <= -'sd4445;
        'd1074: dout <= 'sd445;
        'd1075: dout <= 'sd1284;
        'd1076: dout <= -'sd2749;
        'd1077: dout <= 'sd5324;
        'd1078: dout <= 'sd757;
        'd1079: dout <= 'sd5334;
        'd1080: dout <= 'sd3473;
        'd1081: dout <= -'sd3357;
        'd1082: dout <= 'sd5692;
        'd1083: dout <= 'sd5148;
        'd1084: dout <= -'sd3702;
        'd1085: dout <= -'sd6388;
        'd1086: dout <= 'sd6929;
        'd1087: dout <= -'sd2257;
        'd1088: dout <= -'sd6489;
        'd1089: dout <= -'sd4880;
        'd1090: dout <= -'sd3814;
        'd1091: dout <= -'sd1802;
        'd1092: dout <= 'sd4670;
        'd1093: dout <= 'sd7248;
        'd1094: dout <= 'sd3039;
        'd1095: dout <= 'sd6990;
        'd1096: dout <= -'sd3668;
        'd1097: dout <= -'sd3419;
        'd1098: dout <= 'sd3993;
        'd1099: dout <= -'sd5659;
        'd1100: dout <= -'sd4103;
        'd1101: dout <= -'sd4818;
        'd1102: dout <= 'sd2837;
        'd1103: dout <= 'sd7542;
        'd1104: dout <= -'sd4894;
        'd1105: dout <= -'sd516;
        'd1106: dout <= 'sd4907;
        'd1107: dout <= 'sd2881;
        'd1108: dout <= -'sd7369;
        'd1109: dout <= -'sd4458;
        'd1110: dout <= 'sd427;
        'd1111: dout <= 'sd3755;
        'd1112: dout <= 'sd5185;
        'd1113: dout <= -'sd6827;
        'd1114: dout <= -'sd5710;
        'd1115: dout <= -'sd704;
        'd1116: dout <= -'sd1585;
        'd1117: dout <= -'sd687;
        'd1118: dout <= 'sd2005;
        'd1119: dout <= -'sd4098;
        'd1120: dout <= 'sd7259;
        'd1121: dout <= -'sd5880;
        'd1122: dout <= -'sd5394;
        'd1123: dout <= -'sd5075;
        'd1124: dout <= -'sd7182;
        'd1125: dout <= -'sd5300;
        'd1126: dout <= 'sd5966;
        'd1127: dout <= 'sd1950;
        'd1128: dout <= -'sd7227;
        'd1129: dout <= -'sd3953;
        'd1130: dout <= -'sd6621;
        'd1131: dout <= -'sd2149;
        'd1132: dout <= 'sd4740;
        'd1133: dout <= 'sd3125;
        'd1134: dout <= 'sd1089;
        'd1135: dout <= 'sd6454;
        'd1136: dout <= -'sd3726;
        'd1137: dout <= 'sd2352;
        'd1138: dout <= 'sd2302;
        'd1139: dout <= 'sd6580;
        'd1140: dout <= -'sd3221;
        'd1141: dout <= -'sd6659;
        'd1142: dout <= 'sd7133;
        'd1143: dout <= -'sd2731;
        'd1144: dout <= 'sd1107;
        'd1145: dout <= 'sd6391;
        'd1146: dout <= -'sd5120;
        'd1147: dout <= 'sd1707;
        'd1148: dout <= 'sd1870;
        'd1149: dout <= -'sd4645;
        'd1150: dout <= 'sd6550;
        'd1151: dout <= -'sd1997;
        'd1152: dout <= 'sd528;
        'd1153: dout <= 'sd6311;
        'd1154: dout <= 'sd5605;
        'd1155: dout <= -'sd2531;
        'd1156: dout <= 'sd4913;
        'd1157: dout <= 'sd2479;
        'd1158: dout <= -'sd1179;
        'd1159: dout <= -'sd7341;
        'd1160: dout <= 'sd1773;
        'd1161: dout <= -'sd658;
        'd1162: dout <= 'sd849;
        'd1163: dout <= -'sd5382;
        'd1164: dout <= -'sd1640;
        'd1165: dout <= -'sd6059;
        'd1166: dout <= -'sd5424;
        'd1167: dout <= -'sd1484;
        'd1168: dout <= 'sd3916;
        'd1169: dout <= -'sd1270;
        'd1170: dout <= -'sd319;
        'd1171: dout <= -'sd661;
        'd1172: dout <= 'sd4859;
        'd1173: dout <= -'sd6937;
        'd1174: dout <= 'sd2018;
        'd1175: dout <= 'sd6019;
        'd1176: dout <= 'sd2607;
        'd1177: dout <= 'sd1537;
        'd1178: dout <= -'sd1697;
        'd1179: dout <= 'sd871;
        'd1180: dout <= 'sd2880;
        'd1181: dout <= -'sd6265;
        'd1182: dout <= 'sd338;
        'd1183: dout <= 'sd2625;
        'd1184: dout <= -'sd3184;
        'd1185: dout <= 'sd106;
        'd1186: dout <= 'sd5191;
        'd1187: dout <= -'sd4841;
        'd1188: dout <= 'sd2954;
        'd1189: dout <= -'sd2138;
        'd1190: dout <= 'sd5179;
        'd1191: dout <= -'sd908;
        'd1192: dout <= -'sd6201;
        'd1193: dout <= -'sd1998;
        'd1194: dout <= 'sd4954;
        'd1195: dout <= -'sd5057;
        'd1196: dout <= -'sd6757;
        'd1197: dout <= 'sd7099;
        'd1198: dout <= -'sd1008;
        'd1199: dout <= -'sd3675;
        'd1200: dout <= -'sd3615;
        'd1201: dout <= -'sd4542;
        'd1202: dout <= -'sd3754;
        'd1203: dout <= 'sd6819;
        'd1204: dout <= -'sd5583;
        'd1205: dout <= -'sd884;
        'd1206: dout <= -'sd2470;
        'd1207: dout <= -'sd1548;
        'd1208: dout <= -'sd4571;
        'd1209: dout <= 'sd2029;
        'd1210: dout <= 'sd5961;
        'd1211: dout <= 'sd7127;
        'd1212: dout <= -'sd3911;
        'd1213: dout <= 'sd1033;
        'd1214: dout <= 'sd1269;
        'd1215: dout <= 'sd1865;
        'd1216: dout <= 'sd3091;
        'd1217: dout <= 'sd128;
        'd1218: dout <= 'sd4193;
        'd1219: dout <= -'sd4283;
        'd1220: dout <= 'sd5406;
        'd1221: dout <= 'sd3034;
        'd1222: dout <= -'sd6268;
        'd1223: dout <= -'sd7195;
        'd1224: dout <= 'sd852;
        'd1225: dout <= -'sd2775;
        'd1226: dout <= 'sd3452;
        'd1227: dout <= 'sd6855;
        'd1228: dout <= -'sd1723;
        'd1229: dout <= -'sd1728;
        'd1230: dout <= -'sd956;
        'd1231: dout <= -'sd4918;
        'd1232: dout <= 'sd1743;
        'd1233: dout <= -'sd5216;
        'd1234: dout <= 'sd4333;
        'd1235: dout <= -'sd2372;
        'd1236: dout <= -'sd5512;
        'd1237: dout <= 'sd6507;
        'd1238: dout <= -'sd7256;
        'd1239: dout <= -'sd3721;
        'd1240: dout <= 'sd510;
        'd1241: dout <= -'sd2349;
        'd1242: dout <= -'sd3622;
        'd1243: dout <= 'sd1424;
        'd1244: dout <= -'sd6893;
        'd1245: dout <= 'sd1298;
        'd1246: dout <= 'sd3585;
        'd1247: dout <= 'sd5732;
        'd1248: dout <= -'sd2191;
        'd1249: dout <= -'sd6179;
        'd1250: dout <= -'sd816;
        'd1251: dout <= 'sd2332;
        'd1252: dout <= 'sd6609;
        'd1253: dout <= 'sd866;
        'd1254: dout <= 'sd1110;
        'd1255: dout <= -'sd6487;
        'd1256: dout <= 'sd5615;
        'd1257: dout <= 'sd5849;
        'd1258: dout <= -'sd3069;
        'd1259: dout <= -'sd5217;
        'd1260: dout <= -'sd3775;
        'd1261: dout <= 'sd4110;
        'd1262: dout <= -'sd5698;
        'd1263: dout <= 'sd3699;
        'd1264: dout <= 'sd1751;
        'd1265: dout <= 'sd5141;
        'd1266: dout <= -'sd3449;
        'd1267: dout <= 'sd2383;
        'd1268: dout <= 'sd1436;
        'd1269: dout <= 'sd3843;
        'd1270: dout <= -'sd7179;
        'd1271: dout <= -'sd1513;
        'd1272: dout <= -'sd4415;
        'd1273: dout <= 'sd4416;
        'd1274: dout <= -'sd2402;
        'd1275: dout <= 'sd5305;
        'd1276: dout <= -'sd858;
        'd1277: dout <= 'sd6117;
        'd1278: dout <= 'sd4663;
        'd1279: dout <= 'sd4896;
        'd1280: dout <= -'sd7489;
        'd1281: dout <= -'sd4297;
        'd1282: dout <= 'sd1956;
        'd1283: dout <= 'sd4548;
        'd1284: dout <= 'sd7597;
        'd1285: dout <= 'sd1195;
        'd1286: dout <= -'sd1626;
        'd1287: dout <= -'sd2366;
        'd1288: dout <= -'sd1056;
        'd1289: dout <= -'sd6430;
        'd1290: dout <= 'sd4869;
        'd1291: dout <= -'sd1602;
        'd1292: dout <= 'sd1708;
        'd1293: dout <= 'sd5604;
        'd1294: dout <= -'sd3438;
        'd1295: dout <= 'sd946;
        'd1296: dout <= 'sd1205;
        'd1297: dout <= -'sd7134;
        'd1298: dout <= -'sd6006;
        'd1299: dout <= 'sd2517;
        'd1300: dout <= 'sd1419;
        'd1301: dout <= 'sd5300;
        'd1302: dout <= -'sd7341;
        'd1303: dout <= 'sd6831;
        'd1304: dout <= -'sd4956;
        'd1305: dout <= 'sd3924;
        'd1306: dout <= -'sd7081;
        'd1307: dout <= -'sd3148;
        'd1308: dout <= 'sd1266;
        'd1309: dout <= 'sd3674;
        'd1310: dout <= -'sd1024;
        'd1311: dout <= 'sd715;
        'd1312: dout <= -'sd2251;
        'd1313: dout <= 'sd7337;
        'd1314: dout <= -'sd1709;
        'd1315: dout <= -'sd6466;
        'd1316: dout <= 'sd4364;
        'd1317: dout <= 'sd2926;
        'd1318: dout <= 'sd2452;
        'd1319: dout <= 'sd5965;
        'd1320: dout <= 'sd1318;
        'd1321: dout <= 'sd6637;
        'd1322: dout <= -'sd5160;
        'd1323: dout <= -'sd2079;
        'd1324: dout <= -'sd6091;
        'd1325: dout <= 'sd5824;
        'd1326: dout <= -'sd4587;
        'd1327: dout <= -'sd6744;
        'd1328: dout <= -'sd5481;
        'd1329: dout <= 'sd3681;
        'd1330: dout <= 'sd6646;
        'd1331: dout <= -'sd6932;
        'd1332: dout <= -'sd482;
        'd1333: dout <= -'sd2930;
        'd1334: dout <= 'sd953;
        'd1335: dout <= -'sd6187;
        'd1336: dout <= -'sd2054;
        'd1337: dout <= 'sd236;
        'd1338: dout <= 'sd2793;
        'd1339: dout <= 'sd4143;
        'd1340: dout <= -'sd6276;
        'd1341: dout <= 'sd1323;
        'd1342: dout <= 'sd1189;
        'd1343: dout <= -'sd6788;
        'd1344: dout <= -'sd30;
        'd1345: dout <= 'sd4693;
        'd1346: dout <= 'sd2553;
        'd1347: dout <= -'sd6103;
        'd1348: dout <= -'sd6016;
        'd1349: dout <= 'sd4306;
        'd1350: dout <= 'sd3562;
        'd1351: dout <= 'sd7387;
        'd1352: dout <= 'sd1763;
        'd1353: dout <= -'sd1649;
        'd1354: dout <= 'sd7161;
        'd1355: dout <= 'sd627;
        'd1356: dout <= 'sd484;
        'd1357: dout <= 'sd106;
        'd1358: dout <= 'sd5989;
        'd1359: dout <= -'sd2796;
        'd1360: dout <= 'sd74;
        'd1361: dout <= 'sd6630;
        'd1362: dout <= 'sd3005;
        'd1363: dout <= -'sd3565;
        'd1364: dout <= -'sd5955;
        'd1365: dout <= 'sd6268;
        'd1366: dout <= -'sd4245;
        'd1367: dout <= 'sd6871;
        'd1368: dout <= -'sd1674;
        'd1369: dout <= -'sd1312;
        'd1370: dout <= 'sd1044;
        'd1371: dout <= 'sd3247;
        'd1372: dout <= 'sd5744;
        'd1373: dout <= -'sd1422;
        'd1374: dout <= 'sd6615;
        'd1375: dout <= 'sd4301;
        'd1376: dout <= -'sd2065;
        'd1377: dout <= -'sd2766;
        'd1378: dout <= 'sd3970;
        'd1379: dout <= -'sd503;
        'd1380: dout <= 'sd1329;
        'd1381: dout <= 'sd2422;
        'd1382: dout <= 'sd7541;
        'd1383: dout <= 'sd2917;
        'd1384: dout <= -'sd944;
        'd1385: dout <= -'sd4049;
        'd1386: dout <= -'sd7220;
        'd1387: dout <= -'sd4642;
        'd1388: dout <= 'sd4814;
        'd1389: dout <= 'sd350;
        'd1390: dout <= 'sd6318;
        'd1391: dout <= -'sd5346;
        'd1392: dout <= -'sd3753;
        'd1393: dout <= 'sd5238;
        'd1394: dout <= 'sd7329;
        'd1395: dout <= 'sd316;
        'd1396: dout <= -'sd1927;
        'd1397: dout <= -'sd7012;
        'd1398: dout <= -'sd5363;
        'd1399: dout <= 'sd120;
        'd1400: dout <= -'sd5461;
        'd1401: dout <= -'sd4239;
        'd1402: dout <= -'sd447;
        'd1403: dout <= 'sd2484;
        'd1404: dout <= 'sd1161;
        'd1405: dout <= -'sd1235;
        'd1406: dout <= 'sd988;
        'd1407: dout <= 'sd6024;
        'd1408: dout <= 'sd7379;
        'd1409: dout <= 'sd3406;
        'd1410: dout <= -'sd7252;
        'd1411: dout <= -'sd48;
        'd1412: dout <= -'sd1653;
        'd1413: dout <= -'sd551;
        'd1414: dout <= 'sd7180;
        'd1415: dout <= -'sd5785;
        'd1416: dout <= -'sd7169;
        'd1417: dout <= -'sd5148;
        'd1418: dout <= -'sd1194;
        'd1419: dout <= -'sd6918;
        'd1420: dout <= 'sd933;
        'd1421: dout <= -'sd199;
        'd1422: dout <= -'sd7180;
        'd1423: dout <= 'sd3439;
        'd1424: dout <= -'sd7222;
        'd1425: dout <= 'sd2800;
        'd1426: dout <= 'sd2994;
        'd1427: dout <= 'sd608;
        'd1428: dout <= -'sd5413;
        'd1429: dout <= -'sd28;
        'd1430: dout <= -'sd359;
        'd1431: dout <= -'sd4260;
        'd1432: dout <= -'sd6388;
        'd1433: dout <= -'sd2116;
        'd1434: dout <= -'sd7452;
        'd1435: dout <= 'sd6310;
        'd1436: dout <= -'sd566;
        'd1437: dout <= -'sd3862;
        'd1438: dout <= 'sd2592;
        'd1439: dout <= -'sd4684;
        'd1440: dout <= -'sd4509;
        'd1441: dout <= -'sd6928;
        'd1442: dout <= -'sd376;
        'd1443: dout <= -'sd5086;
        'd1444: dout <= -'sd1471;
        'd1445: dout <= 'sd2652;
        'd1446: dout <= 'sd657;
        'd1447: dout <= 'sd1810;
        'd1448: dout <= -'sd2735;
        'd1449: dout <= 'sd5386;
        'd1450: dout <= 'sd4893;
        'd1451: dout <= 'sd4224;
        'd1452: dout <= -'sd6219;
        'd1453: dout <= 'sd3126;
        'd1454: dout <= 'sd4970;
        'd1455: dout <= -'sd5665;
        'd1456: dout <= -'sd5468;
        'd1457: dout <= -'sd2213;
        'd1458: dout <= 'sd7022;
        'd1459: dout <= 'sd4682;
        'd1460: dout <= 'sd4076;
        'd1461: dout <= 'sd2694;
        'd1462: dout <= -'sd1169;
        'd1463: dout <= 'sd3967;
        'd1464: dout <= -'sd1506;
        'd1465: dout <= 'sd6064;
        'd1466: dout <= 'sd3228;
        'd1467: dout <= 'sd1783;
        'd1468: dout <= 'sd70;
        'd1469: dout <= -'sd3636;
        'd1470: dout <= -'sd1281;
        'd1471: dout <= -'sd4827;
        'd1472: dout <= -'sd1255;
        'd1473: dout <= 'sd6954;
        'd1474: dout <= 'sd4871;
        'd1475: dout <= 'sd624;
        'd1476: dout <= 'sd2671;
        'd1477: dout <= -'sd4339;
        'd1478: dout <= 'sd5351;
        'd1479: dout <= 'sd1209;
        'd1480: dout <= -'sd363;
        'd1481: dout <= -'sd7140;
        'd1482: dout <= 'sd5381;
        'd1483: dout <= -'sd357;
        'd1484: dout <= -'sd2028;
        'd1485: dout <= 'sd514;
        'd1486: dout <= 'sd2184;
        'd1487: dout <= -'sd5867;
        'd1488: dout <= -'sd2336;
        'd1489: dout <= 'sd5536;
        'd1490: dout <= 'sd6076;
        'd1491: dout <= 'sd3715;
        'd1492: dout <= -'sd4721;
        'd1493: dout <= 'sd3542;
        'd1494: dout <= -'sd4767;
        'd1495: dout <= -'sd2509;
        'd1496: dout <= 'sd7530;
        'd1497: dout <= 'sd4077;
        'd1498: dout <= 'sd3060;
        'd1499: dout <= -'sd7521;
        'd1500: dout <= 'sd2955;
        'd1501: dout <= -'sd2547;
        'd1502: dout <= -'sd5909;
        'd1503: dout <= -'sd2241;
        'd1504: dout <= 'sd7345;
        'd1505: dout <= 'sd2425;
        'd1506: dout <= 'sd5751;
        'd1507: dout <= -'sd1459;
        'd1508: dout <= -'sd7650;
        'd1509: dout <= -'sd2228;
        'd1510: dout <= 'sd6330;
        'd1511: dout <= 'sd3001;
        'd1512: dout <= 'sd4214;
        'd1513: dout <= -'sd6509;
        'd1514: dout <= 'sd198;
        'd1515: dout <= 'sd4046;
        'd1516: dout <= -'sd5609;
        'd1517: dout <= 'sd139;
        'd1518: dout <= -'sd3019;
        'd1519: dout <= -'sd7008;
        'd1520: dout <= -'sd432;
        default: dout <= 'sd0;
      endcase
    end
  end

endmodule

